

fn write();
