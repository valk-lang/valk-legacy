
link_static "uv"
