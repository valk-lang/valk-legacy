
value ABE_BOTTOM (3)
value ABE_LEFT (0)
value ABE_RIGHT (2)
value ABE_TOP (1)
value ABM_ACTIVATE (0x00000006)
value ABM_GETAUTOHIDEBAR (0x00000007)
value ABM_GETAUTOHIDEBAREX (0x0000000b)
value ABM_GETSTATE (0x00000004)
value ABM_GETTASKBARPOS (0x00000005)
value ABM_NEW (0x00000000)
value ABM_QUERYPOS (0x00000002)
value ABM_REMOVE (0x00000001)
value ABM_SETAUTOHIDEBAR (0x00000008)
value ABM_SETAUTOHIDEBAREX (0x0000000c)
value ABM_SETPOS (0x00000003)
value ABM_SETSTATE (0x0000000a)
value ABM_WINDOWPOSCHANGED (0x0000009)
value ABN_FULLSCREENAPP (0x0000002)
value ABN_POSCHANGED (0x0000001)
value ABN_STATECHANGE (0x0000000)
value ABN_WINDOWARRANGE (0x0000003)
value ABORTDOC (2)
value ABOVE_NORMAL_PRIORITY_CLASS (0x00008000)
value ABSOLUTE (1)
value ABS_ALWAYSONTOP (0x0000002)
value ABS_AUTOHIDE (0x0000001)
value ACCESS_ALLOWED_ACE_TYPE ((0x0))
value ACCESS_ALLOWED_CALLBACK_ACE_TYPE ((0x9))
value ACCESS_ALLOWED_CALLBACK_OBJECT_ACE_TYPE ((0xB))
value ACCESS_ALLOWED_COMPOUND_ACE_TYPE ((0x4))
value ACCESS_ALLOWED_OBJECT_ACE_TYPE ((0x5))
value ACCESS_DENIED_ACE_TYPE ((0x1))
value ACCESS_DENIED_CALLBACK_ACE_TYPE ((0xA))
value ACCESS_DENIED_CALLBACK_OBJECT_ACE_TYPE ((0xC))
value ACCESS_DENIED_OBJECT_ACE_TYPE ((0x6))
value ACCESS_FILTER_SECURITY_INFORMATION ((0x00000100L))
value ACCESS_MAX_LEVEL (4)
value ACCESS_MAX_MS_ACE_TYPE ((0x8))
value ACCESS_MAX_MS_OBJECT_ACE_TYPE ((0x8))
value ACCESS_MIN_MS_ACE_TYPE ((0x0))
value ACCESS_MIN_MS_OBJECT_ACE_TYPE ((0x5))
value ACCESS_OBJECT_GUID (0)
value ACCESS_PROPERTY_GUID (2)
value ACCESS_PROPERTY_SET_GUID (1)
value ACCESS_REASON_DATA_MASK (0x0000ffff)
value ACCESS_REASON_EXDATA_MASK (0x7f000000)
value ACCESS_REASON_STAGING_MASK (0x80000000)
value ACCESS_REASON_TYPE_MASK (0x00ff0000)
value ACCESS_SYSTEM_SECURITY ((0x01000000L))
value ACE_INHERITED_OBJECT_TYPE_PRESENT (0x2)
value ACE_OBJECT_TYPE_PRESENT (0x1)
value ACL_REVISION ((2))
value ACL_REVISION_DS ((4))
value ACPI_PPM_HARDWARE_ALL (0xFE)
value ACPI_PPM_SOFTWARE_ALL (0xFC)
value ACPI_PPM_SOFTWARE_ANY (0xFD)
value ACTCTX_FLAG_APPLICATION_NAME_VALID ((0x00000020))
value ACTCTX_FLAG_ASSEMBLY_DIRECTORY_VALID ((0x00000004))
value ACTCTX_FLAG_HMODULE_VALID ((0x00000080))
value ACTCTX_FLAG_LANGID_VALID ((0x00000002))
value ACTCTX_FLAG_PROCESSOR_ARCHITECTURE_VALID ((0x00000001))
value ACTCTX_FLAG_RESOURCE_NAME_VALID ((0x00000008))
value ACTCTX_FLAG_SET_PROCESS_DEFAULT ((0x00000010))
value ACTCTX_FLAG_SOURCE_IS_ASSEMBLYREF ((0x00000040))
value ACTIVATIONCONTEXTINFOCLASS (ACTIVATION_CONTEXT_INFO_CLASS)
value ACTIVATION_CONTEXT_BASIC_INFORMATION_DEFINED (1)
value ACTIVATION_CONTEXT_PATH_TYPE_ASSEMBLYREF ((4))
value ACTIVATION_CONTEXT_PATH_TYPE_NONE ((1))
value ACTIVATION_CONTEXT_PATH_TYPE_URL ((3))
value ACTIVATION_CONTEXT_SECTION_APPLICATION_SETTINGS ((10))
value ACTIVATION_CONTEXT_SECTION_ASSEMBLY_INFORMATION ((1))
value ACTIVATION_CONTEXT_SECTION_CLR_SURROGATES ((9))
value ACTIVATION_CONTEXT_SECTION_COMPATIBILITY_INFO ((11))
value ACTIVATION_CONTEXT_SECTION_COM_INTERFACE_REDIRECTION ((5))
value ACTIVATION_CONTEXT_SECTION_COM_PROGID_REDIRECTION ((7))
value ACTIVATION_CONTEXT_SECTION_COM_SERVER_REDIRECTION ((4))
value ACTIVATION_CONTEXT_SECTION_COM_TYPE_LIBRARY_REDIRECTION ((6))
value ACTIVATION_CONTEXT_SECTION_DLL_REDIRECTION ((2))
value ACTIVATION_CONTEXT_SECTION_GLOBAL_OBJECT_RENAME_TABLE ((8))
value ACTIVATION_CONTEXT_SECTION_WINDOW_CLASS_REDIRECTION ((3))
value ACTIVATION_CONTEXT_SECTION_WINRT_ACTIVATABLE_CLASSES ((12))
value ACTIVEOBJECT_STRONG (0x0)
value ACTIVEOBJECT_WEAK (0x1)
value AC_LINE_BACKUP_POWER (0x02)
value AC_LINE_OFFLINE (0x00)
value AC_LINE_ONLINE (0x01)
value AC_LINE_UNKNOWN (0xFF)
value AC_SRC_ALPHA (0x01)
value AC_SRC_OVER (0x00)
value ADDRESS_TAG_BIT (0x40000000000UI64)
value ADDR_ANY (INADDR_ANY)
value AD_CLOCKWISE (2)
value AD_COUNTERCLOCKWISE (1)
value AF_APPLETALK (16)
value AF_ATM (22)
value AF_BAN (21)
value AF_BTH (32)
value AF_CCITT (10)
value AF_CHAOS (5)
value AF_CLUSTER (24)
value AF_DATAKIT (9)
value AF_DLI (13)
value AF_ECMA (8)
value AF_FIREFOX (19)
value AF_HYLINK (15)
value AF_HYPERV (34)
value AF_ICLFXBM (31)
value AF_IMPLINK (3)
value AF_INET (2)
value AF_IPX (AF_NS)
value AF_IRDA (26)
value AF_ISO (7)
value AF_LAT (14)
value AF_LINK (33)
value AF_MAX (35)
value AF_NETBIOS (17)
value AF_NETDES (28)
value AF_NS (6)
value AF_OSI (AF_ISO)
value AF_PUP (4)
value AF_SNA (11)
value AF_TCNMESSAGE (30)
value AF_TCNPROCESS (29)
value AF_UNIX (1)
value AF_UNSPEC (0)
value AF_VOICEVIEW (18)
value AI_ADDRCONFIG (0x00000400)
value AI_ALL (0x00000100)
value AI_BYPASS_DNS_CACHE (0x00000040)
value AI_CANONNAME (0x00000002)
value AI_DISABLE_IDN_ENCODING (0x00080000)
value AI_DNS_ONLY (0x00000010)
value AI_DNS_RESPONSE_HOSTFILE (0x2)
value AI_DNS_RESPONSE_SECURE (0x1)
value AI_DNS_SERVER_TYPE_DOH (0x2)
value AI_DNS_SERVER_TYPE_UDP (0x1)
value AI_DNS_SERVER_UDP_FALLBACK (0x1)
value AI_EXCLUSIVE_CUSTOM_SERVERS (0x00200000)
value AI_EXTENDED (0x80000000)
value AI_FILESERVER (0x00040000)
value AI_FORCE_CLEAR_TEXT (0x00000020)
value AI_FQDN (0x00020000)
value AI_NON_AUTHORITATIVE (0x00004000)
value AI_NUMERICHOST (0x00000004)
value AI_NUMERICSERV (0x00000008)
value AI_PASSIVE (0x00000001)
value AI_REQUIRE_SECURE (0x20000000)
value AI_RESOLUTION_HANDLE (0x40000000)
value AI_RETURN_PREFERRED_NAMES (0x00010000)
value AI_RETURN_RESPONSE_FLAGS (0x10000000)
value AI_RETURN_TTL (0x00000080)
value AI_SECURE (0x00008000)
value AI_SECURE_WITH_FALLBACK (0x00100000)
value ALERT_SYSTEM_CRITICAL (5)
value ALERT_SYSTEM_ERROR (3)
value ALERT_SYSTEM_INFORMATIONAL (1)
value ALERT_SYSTEM_QUERY (4)
value ALERT_SYSTEM_WARNING (2)
value ALG_CLASS_ANY ((0))
value ALG_SID_AES (17)
value ALG_SID_AGREED_KEY_ANY (3)
value ALG_SID_ANY ((0))
value ALG_SID_CAST (6)
value ALG_SID_CYLINK_MEK (12)
value ALG_SID_DES (1)
value ALG_SID_DESX (4)
value ALG_SID_DH_EPHEM (2)
value ALG_SID_DH_SANDF (1)
value ALG_SID_DSS_ANY (0)
value ALG_SID_DSS_DMS (2)
value ALG_SID_DSS_PKCS (1)
value ALG_SID_ECDH (5)
value ALG_SID_ECDH_EPHEM (6)
value ALG_SID_ECDSA (3)
value ALG_SID_ECMQV (1)
value ALG_SID_EXAMPLE (80)
value ALG_SID_HASH_REPLACE_OWF (11)
value ALG_SID_HMAC (9)
value ALG_SID_IDEA (5)
value ALG_SID_KEA (4)
value ALG_SID_MAC (5)
value ALG_SID_RIPEMD (6)
value ALG_SID_RSA_ANY (0)
value ALG_SID_RSA_ENTRUST (3)
value ALG_SID_RSA_MSATWORK (2)
value ALG_SID_RSA_PGP (4)
value ALG_SID_RSA_PKCS (1)
value ALG_SID_SCHANNEL_ENC_KEY (7)
value ALG_SID_SCHANNEL_MAC_KEY (3)
value ALG_SID_SCHANNEL_MASTER_HASH (2)
value ALG_SID_SEAL (2)
value ALG_SID_SHA (4)
value ALG_SID_SKIPJACK (10)
value ALG_SID_TEK (11)
value ALG_SID_THIRDPARTY_ANY ((0))
value ALG_TYPE_ANY ((0))
value ALL_PROCESSOR_GROUPS (0xffff)
value ALTERNATE (1)
value ALTNUMPAD_BIT (0x04000000)
value ANSI_CHARSET (0)
value ANSI_FIXED_FONT (11)
value ANSI_NULL (((CHAR)0))
value ANSI_VAR_FONT (12)
value ANTIALIASED_QUALITY (4)
value ANYSIZE_ARRAY (1)
value APC_LEVEL (1)
value APD_COPY_ALL_FILES (0x00000004)
value APD_COPY_FROM_DIRECTORY (0x00000010)
value APD_COPY_NEW_FILES (0x00000008)
value APD_STRICT_DOWNGRADE (0x00000002)
value APD_STRICT_UPGRADE (0x00000001)
value APIENTRY (WINAPI)
value APPCLASS_MASK (0x0000000FL)
value APPCLASS_MONITOR (0x00000001L)
value APPCLASS_STANDARD (0x00000000L)
value APPCMD_CLIENTONLY (0x00000010L)
value APPCMD_FILTERINITS (0x00000020L)
value APPCMD_MASK (0x00000FF0L)
value APPCOMMAND_BASS_BOOST (20)
value APPCOMMAND_BASS_DOWN (19)
value APPCOMMAND_BASS_UP (21)
value APPCOMMAND_BROWSER_BACKWARD (1)
value APPCOMMAND_BROWSER_FAVORITES (6)
value APPCOMMAND_BROWSER_FORWARD (2)
value APPCOMMAND_BROWSER_HOME (7)
value APPCOMMAND_BROWSER_REFRESH (3)
value APPCOMMAND_BROWSER_SEARCH (5)
value APPCOMMAND_BROWSER_STOP (4)
value APPCOMMAND_CLOSE (31)
value APPCOMMAND_COPY (36)
value APPCOMMAND_CORRECTION_LIST (45)
value APPCOMMAND_CUT (37)
value APPCOMMAND_DELETE (53)
value APPCOMMAND_DICTATE_OR_COMMAND_CONTROL_TOGGLE (43)
value APPCOMMAND_FIND (28)
value APPCOMMAND_FORWARD_MAIL (40)
value APPCOMMAND_HELP (27)
value APPCOMMAND_LAUNCH_MAIL (15)
value APPCOMMAND_LAUNCH_MEDIA_SELECT (16)
value APPCOMMAND_MEDIA_CHANNEL_DOWN (52)
value APPCOMMAND_MEDIA_CHANNEL_UP (51)
value APPCOMMAND_MEDIA_FAST_FORWARD (49)
value APPCOMMAND_MEDIA_NEXTTRACK (11)
value APPCOMMAND_MEDIA_PAUSE (47)
value APPCOMMAND_MEDIA_PLAY (46)
value APPCOMMAND_MEDIA_PLAY_PAUSE (14)
value APPCOMMAND_MEDIA_PREVIOUSTRACK (12)
value APPCOMMAND_MEDIA_RECORD (48)
value APPCOMMAND_MEDIA_REWIND (50)
value APPCOMMAND_MEDIA_STOP (13)
value APPCOMMAND_MICROPHONE_VOLUME_DOWN (25)
value APPCOMMAND_MICROPHONE_VOLUME_MUTE (24)
value APPCOMMAND_MICROPHONE_VOLUME_UP (26)
value APPCOMMAND_MIC_ON_OFF_TOGGLE (44)
value APPCOMMAND_NEW (29)
value APPCOMMAND_OPEN (30)
value APPCOMMAND_PASTE (38)
value APPCOMMAND_PRINT (33)
value APPCOMMAND_REDO (35)
value APPCOMMAND_REPLY_TO_MAIL (39)
value APPCOMMAND_SAVE (32)
value APPCOMMAND_SEND_MAIL (41)
value APPCOMMAND_SPELL_CHECK (42)
value APPCOMMAND_TREBLE_DOWN (22)
value APPCOMMAND_TREBLE_UP (23)
value APPCOMMAND_UNDO (34)
value APPCOMMAND_VOLUME_DOWN (9)
value APPCOMMAND_VOLUME_MUTE (8)
value APPCOMMAND_VOLUME_UP (10)
value APPIDREGFLAGS_AAA_NO_IMPLICIT_ACTIVATE_AS_IU (0x800)
value APPIDREGFLAGS_ACTIVATE_IUSERVER_INDESKTOP (0x1)
value APPIDREGFLAGS_ISSUE_ACTIVATION_RPC_AT_IDENTIFY (0x4)
value APPIDREGFLAGS_IUSERVER_ACTIVATE_IN_CLIENT_SESSION_ONLY (0x20)
value APPIDREGFLAGS_IUSERVER_SELF_SID_IN_LAUNCH_PERMISSION (0x10)
value APPIDREGFLAGS_IUSERVER_UNMODIFIED_LOGON_TOKEN (0x8)
value APPIDREGFLAGS_SECURE_SERVER_PROCESS_SD_AND_BIND (0x2)
value APPLICATION_ERROR_MASK (0x20000000)
value APPMODEL_ERROR_DYNAMIC_PROPERTY_INVALID (15705)
value APPMODEL_ERROR_DYNAMIC_PROPERTY_READ_FAILED (15704)
value APPMODEL_ERROR_NO_APPLICATION (15703)
value APPMODEL_ERROR_NO_MUTABLE_DIRECTORY (15707)
value APPMODEL_ERROR_NO_PACKAGE (15700)
value APPMODEL_ERROR_PACKAGE_IDENTITY_CORRUPT (15702)
value APPMODEL_ERROR_PACKAGE_NOT_AVAILABLE (15706)
value APPMODEL_ERROR_PACKAGE_RUNTIME_CORRUPT (15701)
value APPX_E_BLOCK_HASH_INVALID (_HRESULT_TYPEDEF_(0x80080207L))
value APPX_E_CORRUPT_CONTENT (_HRESULT_TYPEDEF_(0x80080206L))
value APPX_E_DELTA_APPENDED_PACKAGE_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80080210L))
value APPX_E_DELTA_BASELINE_VERSION_MISMATCH (_HRESULT_TYPEDEF_(0x8008020DL))
value APPX_E_DELTA_PACKAGE_MISSING_FILE (_HRESULT_TYPEDEF_(0x8008020EL))
value APPX_E_DIGEST_MISMATCH (_HRESULT_TYPEDEF_(0x80080219L))
value APPX_E_FILE_COMPRESSION_MISMATCH (_HRESULT_TYPEDEF_(0x80080214L))
value APPX_E_INTERLEAVING_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80080201L))
value APPX_E_INVALID_APPINSTALLER (_HRESULT_TYPEDEF_(0x8008020CL))
value APPX_E_INVALID_BLOCKMAP (_HRESULT_TYPEDEF_(0x80080205L))
value APPX_E_INVALID_CONTENTGROUPMAP (_HRESULT_TYPEDEF_(0x8008020BL))
value APPX_E_INVALID_DELTA_PACKAGE (_HRESULT_TYPEDEF_(0x8008020FL))
value APPX_E_INVALID_ENCRYPTION_EXCLUSION_FILE_LIST (_HRESULT_TYPEDEF_(0x80080216L))
value APPX_E_INVALID_KEY_INFO (_HRESULT_TYPEDEF_(0x8008020AL))
value APPX_E_INVALID_MANIFEST (_HRESULT_TYPEDEF_(0x80080204L))
value APPX_E_INVALID_PACKAGESIGNCONFIG (_HRESULT_TYPEDEF_(0x80080212L))
value APPX_E_INVALID_PACKAGE_FOLDER_ACLS (_HRESULT_TYPEDEF_(0x80080217L))
value APPX_E_INVALID_PACKAGING_LAYOUT (_HRESULT_TYPEDEF_(0x80080211L))
value APPX_E_INVALID_PAYLOAD_PACKAGE_EXTENSION (_HRESULT_TYPEDEF_(0x80080215L))
value APPX_E_INVALID_PUBLISHER_BRIDGING (_HRESULT_TYPEDEF_(0x80080218L))
value APPX_E_INVALID_SIP_CLIENT_DATA (_HRESULT_TYPEDEF_(0x80080209L))
value APPX_E_MISSING_REQUIRED_FILE (_HRESULT_TYPEDEF_(0x80080203L))
value APPX_E_PACKAGING_INTERNAL (_HRESULT_TYPEDEF_(0x80080200L))
value APPX_E_RELATIONSHIPS_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80080202L))
value APPX_E_REQUESTED_RANGE_TOO_LARGE (_HRESULT_TYPEDEF_(0x80080208L))
value APPX_E_RESOURCESPRI_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80080213L))
value APP_LOCAL_DEVICE_ID_SIZE (32)
value ARABIC_CHARSET (178)
value ARM_CACHE_ALIGNMENT_SIZE (128)
value ARW_BOTTOMLEFT (0x0000L)
value ARW_BOTTOMRIGHT (0x0001L)
value ARW_DOWN (0x0004L)
value ARW_HIDE (0x0008L)
value ARW_LEFT (0x0000L)
value ARW_RIGHT (0x0000L)
value ARW_STARTMASK (0x0003L)
value ARW_STARTRIGHT (0x0001L)
value ARW_STARTTOP (0x0002L)
value ARW_TOPLEFT (0x0002L)
value ARW_TOPRIGHT (0x0003L)
value ARW_UP (0x0004L)
value ASFW_ANY (((DWORD)-1))
value ASPECTX (40)
value ASPECTXY (44)
value ASPECTY (42)
value ASPECT_FILTERING (0x0001)
value ASSEMBLY_DLL_REDIRECTION_DETAILED_INFORMATION (ASSEMBLY_FILE_DETAILED_INFORMATION)
value ASSERT_ALTERNATE (0x9)
value ASSERT_PRIMARY (0x8)
value ASYNCH (0x80)
value ASYNC_MODE_COMPATIBILITY (0x00000001L)
value ASYNC_MODE_DEFAULT (0x00000000L)
value ATAPI_ID_CMD (0xA1)
value ATF_ONOFFFEEDBACK (0x00000002)
value ATF_TIMEOUTON (0x00000001)
value ATOM_FLAG_GLOBAL (0x2)
value ATTACH_PARENT_PROCESS (((DWORD)-1))
value ATTRIBUTE_SECURITY_INFORMATION ((0x00000020L))
value ATTR_CONVERTED (0x02)
value ATTR_FIXEDCONVERTED (0x05)
value ATTR_INPUT (0x00)
value ATTR_INPUT_ERROR (0x04)
value ATTR_TARGET_CONVERTED (0x01)
value ATTR_TARGET_NOTCONVERTED (0x03)
value AT_KEYEXCHANGE (1)
value AT_SIGNATURE (2)
value AUDIT_ALLOW_NO_PRIVILEGE (0x1)
value AUTHTYPE_CLIENT (1)
value AUTHTYPE_SERVER (2)
value AUXCAPS_AUXIN (2)
value AUXCAPS_CDAUDIO (1)
value AUXCAPS_LRVOLUME (0x0002)
value AUXCAPS_VOLUME (0x0001)
value AUX_MAPPER (((UINT)-1))
value AW_ACTIVATE (0x00020000)
value AW_BLEND (0x00080000)
value AW_CENTER (0x00000010)
value AW_HIDE (0x00010000)
value AW_HOR_NEGATIVE (0x00000002)
value AW_HOR_POSITIVE (0x00000001)
value AW_SLIDE (0x00040000)
value AW_VER_NEGATIVE (0x00000008)
value AW_VER_POSITIVE (0x00000004)
value BACKGROUND_BLUE (0x0010)
value BACKGROUND_GREEN (0x0020)
value BACKGROUND_INTENSITY (0x0080)
value BACKGROUND_RED (0x0040)
value BACKUP_ALTERNATE_DATA (0x00000004)
value BACKUP_DATA (0x00000001)
value BACKUP_EA_DATA (0x00000002)
value BACKUP_GHOSTED_FILE_EXTENTS (0x0000000b)
value BACKUP_INVALID (0x00000000)
value BACKUP_LINK (0x00000005)
value BACKUP_OBJECT_ID (0x00000007)
value BACKUP_PROPERTY_DATA (0x00000006)
value BACKUP_REPARSE_DATA (0x00000008)
value BACKUP_SECURITY_DATA (0x00000003)
value BACKUP_SECURITY_INFORMATION ((0x00010000L))
value BACKUP_SPARSE_BLOCK (0x00000009)
value BACKUP_TXFS_DATA (0x0000000a)
value BALTIC_CHARSET (186)
value BANDINFO (24)
value BASE_PROTOCOL (1)
value BASE_SEARCH_PATH_DISABLE_SAFE_SEARCHMODE (0x10000)
value BASE_SEARCH_PATH_ENABLE_SAFE_SEARCHMODE (0x1)
value BASE_SEARCH_PATH_PERMANENT (0x8000)
value BASIC_CONSTRAINTS_CERT_CHAIN_POLICY_CA_FLAG (0x80000000)
value BASIC_CONSTRAINTS_CERT_CHAIN_POLICY_END_ENTITY_FLAG (0x40000000)
value BATTERY_DISCHARGE_FLAGS_ENABLE (0x80000000)
value BATTERY_DISCHARGE_FLAGS_EVENTCODE_MASK (0x00000007)
value BATTERY_FLAG_CHARGING (0x08)
value BATTERY_FLAG_CRITICAL (0x04)
value BATTERY_FLAG_HIGH (0x01)
value BATTERY_FLAG_LOW (0x02)
value BATTERY_FLAG_NO_BATTERY (0x80)
value BATTERY_FLAG_UNKNOWN (0xFF)
value BATTERY_LIFE_UNKNOWN (0xFFFFFFFF)
value BATTERY_PERCENTAGE_UNKNOWN (0xFF)
value BAUD_USER (((DWORD)0x10000000))
value BCRYPTBUFFER_VERSION (0)
value BCRYPT_AES_CMAC_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000101))
value BCRYPT_AES_GMAC_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000111))
value BCRYPT_ALG_HANDLE_HMAC_FLAG (0x00000008)
value BCRYPT_ASYMMETRIC_ENCRYPTION_INTERFACE (0x00000003)
value BCRYPT_ASYMMETRIC_ENCRYPTION_OPERATION (0x00000004)
value BCRYPT_AUTHENTICATED_CIPHER_MODE_INFO_VERSION (1)
value BCRYPT_AUTH_MODE_CHAIN_CALLS_FLAG (0x00000001)
value BCRYPT_AUTH_MODE_IN_PROGRESS_FLAG (0x00000002)
value BCRYPT_BLOCK_PADDING (0x00000001)
value BCRYPT_BUFFERS_LOCKED_FLAG (0x00000040)
value BCRYPT_CAPI_AES_FLAG (0x00000010)
value BCRYPT_CAPI_KDF_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000321))
value BCRYPT_CIPHER_INTERFACE (0x00000001)
value BCRYPT_CIPHER_OPERATION (0x00000001)
value BCRYPT_DESX_CBC_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000221))
value BCRYPT_DESX_CFB_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000241))
value BCRYPT_DESX_ECB_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000231))
value BCRYPT_DES_CFB_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000211))
value BCRYPT_DES_ECB_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000201))
value BCRYPT_DH_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000281))
value BCRYPT_DH_PARAMETERS_MAGIC (0x4d504844)
value BCRYPT_DH_PRIVATE_MAGIC (0x56504844)
value BCRYPT_DH_PUBLIC_MAGIC (0x42504844)
value BCRYPT_DSA_PARAMETERS_MAGIC (0x4d505344)
value BCRYPT_DSA_PRIVATE_MAGIC (0x56505344)
value BCRYPT_DSA_PUBLIC_MAGIC (0x42505344)
value BCRYPT_ECC_PARAMETERS_MAGIC (0x50434345)
value BCRYPT_ECDH_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000291))
value BCRYPT_ECDH_PRIVATE_GENERIC_MAGIC (0x564B4345)
value BCRYPT_ECDH_PUBLIC_GENERIC_MAGIC (0x504B4345)
value BCRYPT_ECDSA_PRIVATE_GENERIC_MAGIC (0x56444345)
value BCRYPT_ECDSA_PUBLIC_GENERIC_MAGIC (0x50444345)
value BCRYPT_ENABLE_INCOMPATIBLE_FIPS_CHECKS (0x00000100)
value BCRYPT_EXTENDED_KEYSIZE (0x00000080)
value BCRYPT_GENERATE_IV (0x00000020)
value BCRYPT_HASH_INTERFACE (0x00000002)
value BCRYPT_HASH_OPERATION (0x00000002)
value BCRYPT_HASH_REUSABLE_FLAG (0x00000020)
value BCRYPT_HKDF_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000391))
value BCRYPT_KEY_DATA_BLOB_MAGIC (0x4d42444b)
value BCRYPT_KEY_DERIVATION_INTERFACE (0x00000007)
value BCRYPT_KEY_DERIVATION_OPERATION (0x00000040)
value BCRYPT_KEY_VALIDATION_RANGE (0x00000010)
value BCRYPT_KEY_VALIDATION_RANGE_AND_ORDER (0x00000018)
value BCRYPT_KEY_VALIDATION_REGENERATE (0x00000020)
value BCRYPT_MULTI_FLAG (0x00000040)
value BCRYPT_NO_KEY_VALIDATION (0x00000008)
value BCRYPT_OBJECT_ALIGNMENT (16)
value BCRYPT_PAD_NONE (0x00000001)
value BCRYPT_PAD_OAEP (0x00000004)
value BCRYPT_PAD_PSS (0x00000008)
value BCRYPT_PRIVATE_KEY_FLAG (0x00000002)
value BCRYPT_PROV_DISPATCH (0x00000001)
value BCRYPT_PUBLIC_KEY_FLAG (0x00000001)
value BCRYPT_RNG_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000081))
value BCRYPT_RNG_INTERFACE (0x00000006)
value BCRYPT_RNG_OPERATION (0x00000020)
value BCRYPT_RNG_USE_ENTROPY_IN_BUFFER (0x00000001)
value BCRYPT_RSAFULLPRIVATE_MAGIC (0x33415352)
value BCRYPT_RSAPRIVATE_MAGIC (0x32415352)
value BCRYPT_RSAPUBLIC_MAGIC (0x31415352)
value BCRYPT_RSA_SIGN_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000311))
value BCRYPT_SECRET_AGREEMENT_INTERFACE (0x00000004)
value BCRYPT_SECRET_AGREEMENT_OPERATION (0x00000008)
value BCRYPT_SIGNATURE_INTERFACE (0x00000005)
value BCRYPT_SIGNATURE_OPERATION (0x00000010)
value BCRYPT_SUPPORTED_PAD_OAEP (0x00000008)
value BCRYPT_SUPPORTED_PAD_PSS (0x00000010)
value BCRYPT_SUPPORTED_PAD_ROUTER (0x00000001)
value BCRYPT_TLS_CBC_HMAC_VERIFY_FLAG (0x00000004)
value BCRYPT_USE_SYSTEM_PREFERRED_RNG (0x00000002)
value BCRYPT_XTS_AES_ALG_HANDLE (((BCRYPT_ALG_HANDLE) 0x00000381))
value BDR_INNER ((BDR_RAISEDINNER | BDR_SUNKENINNER))
value BDR_OUTER ((BDR_RAISEDOUTER | BDR_SUNKENOUTER))
value BDR_RAISED ((BDR_RAISEDOUTER | BDR_RAISEDINNER))
value BDR_RAISEDINNER (0x0004)
value BDR_RAISEDOUTER (0x0001)
value BDR_SUNKEN ((BDR_SUNKENOUTER | BDR_SUNKENINNER))
value BDR_SUNKENINNER (0x0008)
value BDR_SUNKENOUTER (0x0002)
value BEGIN_PATH (4096)
value BELOW_NORMAL_PRIORITY_CLASS (0x00004000)
value BF_ADJUST (0x2000)
value BF_BOTTOM (0x0008)
value BF_BOTTOMLEFT ((BF_BOTTOM | BF_LEFT))
value BF_BOTTOMRIGHT ((BF_BOTTOM | BF_RIGHT))
value BF_DIAGONAL (0x0010)
value BF_DIAGONAL_ENDBOTTOMLEFT ((BF_DIAGONAL | BF_BOTTOM | BF_LEFT))
value BF_DIAGONAL_ENDBOTTOMRIGHT ((BF_DIAGONAL | BF_BOTTOM | BF_RIGHT))
value BF_DIAGONAL_ENDTOPLEFT ((BF_DIAGONAL | BF_TOP | BF_LEFT))
value BF_DIAGONAL_ENDTOPRIGHT ((BF_DIAGONAL | BF_TOP | BF_RIGHT))
value BF_FLAT (0x4000)
value BF_LEFT (0x0001)
value BF_MIDDLE (0x0800)
value BF_MONO (0x8000)
value BF_RECT ((BF_LEFT | BF_TOP | BF_RIGHT | BF_BOTTOM))
value BF_RIGHT (0x0004)
value BF_SOFT (0x1000)
value BF_TOP (0x0002)
value BF_TOPLEFT ((BF_TOP | BF_LEFT))
value BF_TOPRIGHT ((BF_TOP | BF_RIGHT))
value BIDI_ACCESS_ADMINISTRATOR (0x1)
value BIDI_ACCESS_USER (0x2)
value BIGENDIAN (0x0000)
value BINDF_DONTPUTINCACHE (32)
value BINDF_DONTUSECACHE (16)
value BINDF_NOCOPYDATA (128)
value BITSPIXEL (12)
value BI_BITFIELDS (3)
value BI_JPEG (4)
value BI_PNG (5)
value BI_RGB (0)
value BKMODE_LAST (2)
value BLACKNESS ((DWORD)0x00000042)
value BLACKONWHITE (1)
value BLACK_BRUSH (4)
value BLACK_PEN (7)
value BLTALIGNMENT (119)
value BM_CLICK (0x00F5)
value BM_GETCHECK (0x00F0)
value BM_GETIMAGE (0x00F6)
value BM_GETSTATE (0x00F2)
value BM_SETCHECK (0x00F1)
value BM_SETDONTCLICK (0x00F8)
value BM_SETIMAGE (0x00F7)
value BM_SETSTATE (0x00F3)
value BM_SETSTYLE (0x00F4)
value BN_CLICKED (0)
value BN_DBLCLK (BN_DOUBLECLICKED)
value BN_DISABLE (4)
value BN_DOUBLECLICKED (5)
value BN_HILITE (2)
value BN_KILLFOCUS (7)
value BN_PAINT (1)
value BN_PUSHED (BN_HILITE)
value BN_SETFOCUS (6)
value BN_UNHILITE (3)
value BN_UNPUSHED (BN_UNHILITE)
value BOLD_FONTTYPE (0x0100)
value BROADCAST_QUERY_DENY (0x424D5144)
value BSF_ALLOWSFW (0x00000080)
value BSF_FLUSHDISK (0x00000004)
value BSF_FORCEIFHUNG (0x00000020)
value BSF_IGNORECURRENTTASK (0x00000002)
value BSF_LUID (0x00000400)
value BSF_NOHANG (0x00000008)
value BSF_NOTIMEOUTIFNOTHUNG (0x00000040)
value BSF_POSTMESSAGE (0x00000010)
value BSF_QUERY (0x00000001)
value BSF_RETURNHDESK (0x00000200)
value BSF_SENDNOTIFYMESSAGE (0x00000100)
value BSM_ALLCOMPONENTS (0x00000000)
value BSM_ALLDESKTOPS (0x00000010)
value BSM_APPLICATIONS (0x00000008)
value BSM_INSTALLABLEDRIVERS (0x00000004)
value BSM_NETDRIVER (0x00000002)
value BSM_VXDS (0x00000001)
value BST_CHECKED (0x0001)
value BST_FOCUS (0x0008)
value BST_INDETERMINATE (0x0002)
value BST_PUSHED (0x0004)
value BST_UNCHECKED (0x0000)
value BS_AUTOCHECKBOX (0x00000003L)
value BS_AUTORADIOBUTTON (0x00000009L)
value BS_BITMAP (0x00000080L)
value BS_BOTTOM (0x00000800L)
value BS_CENTER (0x00000300L)
value BS_CHECKBOX (0x00000002L)
value BS_DEFPUSHBUTTON (0x00000001L)
value BS_DIBPATTERN (5)
value BS_DIBPATTERNPT (6)
value BS_FLAT (0x00008000L)
value BS_GROUPBOX (0x00000007L)
value BS_HATCHED (2)
value BS_HOLLOW (BS_NULL)
value BS_ICON (0x00000040L)
value BS_INDEXED (4)
value BS_LEFT (0x00000100L)
value BS_LEFTTEXT (0x00000020L)
value BS_MONOPATTERN (9)
value BS_MULTILINE (0x00002000L)
value BS_NOTIFY (0x00004000L)
value BS_NULL (1)
value BS_OWNERDRAW (0x0000000BL)
value BS_PATTERN (3)
value BS_PUSHBOX (0x0000000AL)
value BS_PUSHBUTTON (0x00000000L)
value BS_PUSHLIKE (0x00001000L)
value BS_RADIOBUTTON (0x00000004L)
value BS_RIGHT (0x00000200L)
value BS_RIGHTBUTTON (BS_LEFTTEXT)
value BS_SOLID (0)
value BS_TEXT (0x00000000L)
value BS_TOP (0x00000400L)
value BS_TYPEMASK (0x0000000FL)
value BS_USERBUTTON (0x00000008L)
value BS_VCENTER (0x00000C00L)
value BT_E_SPURIOUS_ACTIVATION (_HRESULT_TYPEDEF_(0x80080300L))
value BUFSIZ (512)
value CACHE_E_FIRST (0x80040170L)
value CACHE_E_LAST (0x8004017FL)
value CACHE_E_NOCACHE_UPDATED (_HRESULT_TYPEDEF_(0x80040170L))
value CACHE_FULLY_ASSOCIATIVE (0xFF)
value CACHE_S_FIRST (0x00040170L)
value CACHE_S_FORMATETC_NOTSUPPORTED (_HRESULT_TYPEDEF_(0x00040170L))
value CACHE_S_LAST (0x0004017FL)
value CACHE_S_SAMECACHE (_HRESULT_TYPEDEF_(0x00040171L))
value CACHE_S_SOMECACHES_NOTUPDATED (_HRESULT_TYPEDEF_(0x00040172L))
value CADV_LATEACK (0xFFFF)
value CALERT_SYSTEM (6)
value CALG_AES ((ALG_CLASS_DATA_ENCRYPT|ALG_TYPE_BLOCK|ALG_SID_AES))
value CALG_AGREEDKEY_ANY ((ALG_CLASS_KEY_EXCHANGE|ALG_TYPE_DH|ALG_SID_AGREED_KEY_ANY))
value CALG_CYLINK_MEK ((ALG_CLASS_DATA_ENCRYPT|ALG_TYPE_BLOCK|ALG_SID_CYLINK_MEK))
value CALG_DES ((ALG_CLASS_DATA_ENCRYPT|ALG_TYPE_BLOCK|ALG_SID_DES))
value CALG_DESX ((ALG_CLASS_DATA_ENCRYPT|ALG_TYPE_BLOCK|ALG_SID_DESX))
value CALG_DH_EPHEM ((ALG_CLASS_KEY_EXCHANGE|ALG_TYPE_DH|ALG_SID_DH_EPHEM))
value CALG_DH_SF ((ALG_CLASS_KEY_EXCHANGE|ALG_TYPE_DH|ALG_SID_DH_SANDF))
value CALG_DSS_SIGN ((ALG_CLASS_SIGNATURE | ALG_TYPE_DSS | ALG_SID_DSS_ANY))
value CALG_ECDH ((ALG_CLASS_KEY_EXCHANGE | ALG_TYPE_DH | ALG_SID_ECDH))
value CALG_ECDH_EPHEM ((ALG_CLASS_KEY_EXCHANGE | ALG_TYPE_ECDH | ALG_SID_ECDH_EPHEM))
value CALG_ECDSA ((ALG_CLASS_SIGNATURE | ALG_TYPE_DSS | ALG_SID_ECDSA))
value CALG_ECMQV ((ALG_CLASS_KEY_EXCHANGE | ALG_TYPE_ANY | ALG_SID_ECMQV))
value CALG_HASH_REPLACE_OWF ((ALG_CLASS_HASH | ALG_TYPE_ANY | ALG_SID_HASH_REPLACE_OWF))
value CALG_HMAC ((ALG_CLASS_HASH | ALG_TYPE_ANY | ALG_SID_HMAC))
value CALG_KEA_KEYX ((ALG_CLASS_KEY_EXCHANGE|ALG_TYPE_DH|ALG_SID_KEA))
value CALG_MAC ((ALG_CLASS_HASH | ALG_TYPE_ANY | ALG_SID_MAC))
value CALG_NO_SIGN ((ALG_CLASS_SIGNATURE | ALG_TYPE_ANY | ALG_SID_ANY))
value CALG_NULLCIPHER ((ALG_CLASS_DATA_ENCRYPT | ALG_TYPE_ANY | 0))
value CALG_OID_INFO_CNG_ONLY (0xFFFFFFFF)
value CALG_OID_INFO_PARAMETERS (0xFFFFFFFE)
value CALG_RSA_KEYX ((ALG_CLASS_KEY_EXCHANGE|ALG_TYPE_RSA|ALG_SID_RSA_ANY))
value CALG_RSA_SIGN ((ALG_CLASS_SIGNATURE | ALG_TYPE_RSA | ALG_SID_RSA_ANY))
value CALG_SCHANNEL_ENC_KEY ((ALG_CLASS_MSG_ENCRYPT|ALG_TYPE_SECURECHANNEL|ALG_SID_SCHANNEL_ENC_KEY))
value CALG_SCHANNEL_MAC_KEY ((ALG_CLASS_MSG_ENCRYPT|ALG_TYPE_SECURECHANNEL|ALG_SID_SCHANNEL_MAC_KEY))
value CALG_SCHANNEL_MASTER_HASH ((ALG_CLASS_MSG_ENCRYPT|ALG_TYPE_SECURECHANNEL|ALG_SID_SCHANNEL_MASTER_HASH))
value CALG_SEAL ((ALG_CLASS_DATA_ENCRYPT|ALG_TYPE_STREAM|ALG_SID_SEAL))
value CALG_SHA ((ALG_CLASS_HASH | ALG_TYPE_ANY | ALG_SID_SHA))
value CALG_SKIPJACK ((ALG_CLASS_DATA_ENCRYPT|ALG_TYPE_BLOCK|ALG_SID_SKIPJACK))
value CALG_TEK ((ALG_CLASS_DATA_ENCRYPT|ALG_TYPE_BLOCK|ALG_SID_TEK))
value CALG_THIRDPARTY_CIPHER ((ALG_CLASS_DATA_ENCRYPT | ALG_TYPE_THIRDPARTY | ALG_SID_THIRDPARTY_ANY))
value CALG_THIRDPARTY_HASH ((ALG_CLASS_HASH | ALG_TYPE_THIRDPARTY | ALG_SID_THIRDPARTY_ANY))
value CALG_THIRDPARTY_KEY_EXCHANGE ((ALG_CLASS_KEY_EXCHANGE | ALG_TYPE_THIRDPARTY | ALG_SID_THIRDPARTY_ANY))
value CALG_THIRDPARTY_SIGNATURE ((ALG_CLASS_SIGNATURE | ALG_TYPE_THIRDPARTY | ALG_SID_THIRDPARTY_ANY))
value CALINFO_ENUMPROC (CALINFO_ENUMPROCA)
value CALINFO_ENUMPROCEX (CALINFO_ENUMPROCEXA)
value CALLBACK_CHUNK_FINISHED (0x00000000)
value CALLBACK_STREAM_SWITCH (0x00000001)
value CALLBACK_THREAD ((CALLBACK_TASK))
value CALL_PENDING (0x02)
value CAL_GREGORIAN (1)
value CAL_GREGORIAN_ARABIC (10)
value CAL_GREGORIAN_ME_FRENCH (9)
value CAL_GREGORIAN_US (2)
value CAL_GREGORIAN_XLIT_ENGLISH (11)
value CAL_GREGORIAN_XLIT_FRENCH (12)
value CAL_HEBREW (8)
value CAL_HIJRI (6)
value CAL_ICALINTVALUE (0x00000001)
value CAL_ITWODIGITYEARMAX (0x00000030)
value CAL_IYEAROFFSETRANGE (0x00000003)
value CAL_JAPAN (3)
value CAL_KOREA (5)
value CAL_NOUSEROVERRIDE (LOCALE_NOUSEROVERRIDE)
value CAL_PERSIAN (22)
value CAL_RETURN_GENITIVE_NAMES (LOCALE_RETURN_GENITIVE_NAMES)
value CAL_RETURN_NUMBER (LOCALE_RETURN_NUMBER)
value CAL_SABBREVERASTRING (0x00000039)
value CAL_SCALNAME (0x00000002)
value CAL_SENGLISHABBREVERANAME (0x0000003c)
value CAL_SENGLISHERANAME (0x0000003b)
value CAL_SERASTRING (0x00000004)
value CAL_SJAPANESEERAFIRSTYEAR (0x0000003d)
value CAL_SLONGDATE (0x00000006)
value CAL_SMONTHDAY (0x00000038)
value CAL_SRELATIVELONGDATE (0x0000003a)
value CAL_SSHORTDATE (0x00000005)
value CAL_SYEARMONTH (0x0000002f)
value CAL_TAIWAN (4)
value CAL_THAI (7)
value CAL_UMALQURA (23)
value CAL_USE_CP_ACP (LOCALE_USE_CP_ACP)
value CAPSLOCK_ON (0x0080)
value CAPTUREBLT ((DWORD)0x40000000)
value CAP_ATAPI_ID_CMD (2)
value CAP_ATA_ID_CMD (1)
value CAP_SMART_CMD (4)
value CAT_E_CATIDNOEXIST (_HRESULT_TYPEDEF_(0x80040160L))
value CAT_E_FIRST (0x80040160L)
value CAT_E_LAST (0x80040161L)
value CAT_E_NODESCRIPTION (_HRESULT_TYPEDEF_(0x80040161L))
value CA_LOG_FILTER (0x0002)
value CA_NEGATIVE (0x0001)
value CBF_FAIL_ADVISES (0x00004000)
value CBF_FAIL_ALLSVRXACTIONS (0x0003f000)
value CBF_FAIL_CONNECTIONS (0x00002000)
value CBF_FAIL_EXECUTES (0x00008000)
value CBF_FAIL_POKES (0x00010000)
value CBF_FAIL_REQUESTS (0x00020000)
value CBF_FAIL_SELFCONNECTIONS (0x00001000)
value CBF_SKIP_ALLNOTIFICATIONS (0x003c0000)
value CBF_SKIP_CONNECT_CONFIRMS (0x00040000)
value CBF_SKIP_DISCONNECTS (0x00200000)
value CBF_SKIP_REGISTRATIONS (0x00080000)
value CBF_SKIP_UNREGISTRATIONS (0x00100000)
value CBM_INIT (0x04L)
value CBN_CLOSEUP (8)
value CBN_DBLCLK (2)
value CBN_DROPDOWN (7)
value CBN_EDITCHANGE (5)
value CBN_EDITUPDATE (6)
value CBN_ERRSPACE ((-1))
value CBN_KILLFOCUS (4)
value CBN_SELCHANGE (1)
value CBN_SELENDCANCEL (10)
value CBN_SELENDOK (9)
value CBN_SETFOCUS (3)
value CBR_BLOCK (((HDDEDATA)-1))
value CBS_AUTOHSCROLL (0x0040L)
value CBS_DISABLENOSCROLL (0x0800L)
value CBS_DROPDOWN (0x0002L)
value CBS_DROPDOWNLIST (0x0003L)
value CBS_HASSTRINGS (0x0200L)
value CBS_LOWERCASE (0x4000L)
value CBS_NOINTEGRALHEIGHT (0x0400L)
value CBS_OEMCONVERT (0x0080L)
value CBS_OWNERDRAWFIXED (0x0010L)
value CBS_OWNERDRAWVARIABLE (0x0020L)
value CBS_SIMPLE (0x0001L)
value CBS_SORT (0x0100L)
value CBS_UPPERCASE (0x2000L)
value CB_ADDSTRING (0x0143)
value CB_DELETESTRING (0x0144)
value CB_DIR (0x0145)
value CB_ERR ((-1))
value CB_ERRSPACE ((-2))
value CB_FINDSTRING (0x014C)
value CB_FINDSTRINGEXACT (0x0158)
value CB_GETCOMBOBOXINFO (0x0164)
value CB_GETCOUNT (0x0146)
value CB_GETCURSEL (0x0147)
value CB_GETDROPPEDCONTROLRECT (0x0152)
value CB_GETDROPPEDSTATE (0x0157)
value CB_GETDROPPEDWIDTH (0x015f)
value CB_GETEDITSEL (0x0140)
value CB_GETEXTENDEDUI (0x0156)
value CB_GETHORIZONTALEXTENT (0x015d)
value CB_GETITEMDATA (0x0150)
value CB_GETITEMHEIGHT (0x0154)
value CB_GETLBTEXT (0x0148)
value CB_GETLBTEXTLEN (0x0149)
value CB_GETLOCALE (0x015A)
value CB_GETTOPINDEX (0x015b)
value CB_INITSTORAGE (0x0161)
value CB_INSERTSTRING (0x014A)
value CB_LIMITTEXT (0x0141)
value CB_MSGMAX (0x0165)
value CB_OKAY (0)
value CB_RESETCONTENT (0x014B)
value CB_SELECTSTRING (0x014D)
value CB_SETCURSEL (0x014E)
value CB_SETDROPPEDWIDTH (0x0160)
value CB_SETEDITSEL (0x0142)
value CB_SETEXTENDEDUI (0x0155)
value CB_SETHORIZONTALEXTENT (0x015e)
value CB_SETITEMDATA (0x0151)
value CB_SETITEMHEIGHT (0x0153)
value CB_SETLOCALE (0x0159)
value CB_SETTOPINDEX (0x015c)
value CB_SHOWDROPDOWN (0x014F)
value CCERR_CHOOSECOLORCODES (0x5000)
value CCHDEVICENAME (32)
value CCHFORMNAME (32)
value CCHILDREN_SCROLLBAR (5)
value CCHILDREN_TITLEBAR (5)
value CCH_MAX_PROPSTG_NAME (31)
value CC_ANYCOLOR (0x00000100)
value CC_CHORD (4)
value CC_CIRCLES (1)
value CC_ELLIPSES (8)
value CC_ENABLEHOOK (0x00000010)
value CC_ENABLETEMPLATE (0x00000020)
value CC_ENABLETEMPLATEHANDLE (0x00000040)
value CC_FULLOPEN (0x00000002)
value CC_INTERIORS (128)
value CC_NONE (0)
value CC_PIE (2)
value CC_PREVENTFULLOPEN (0x00000004)
value CC_RGBINIT (0x00000001)
value CC_ROUNDRECT (256)
value CC_SHOWHELP (0x00000008)
value CC_SOLIDCOLOR (0x00000080)
value CC_STYLED (32)
value CC_WIDE (16)
value CC_WIDESTYLED (64)
value CDB_SIZE (16)
value CDERR_DIALOGFAILURE (0xFFFF)
value CDERR_FINDRESFAILURE (0x0006)
value CDERR_GENERALCODES (0x0000)
value CDERR_INITIALIZATION (0x0002)
value CDERR_LOADRESFAILURE (0x0007)
value CDERR_LOADSTRFAILURE (0x0005)
value CDERR_LOCKRESFAILURE (0x0008)
value CDERR_MEMALLOCFAILURE (0x0009)
value CDERR_MEMLOCKFAILURE (0x000A)
value CDERR_NOHINSTANCE (0x0004)
value CDERR_NOHOOK (0x000B)
value CDERR_NOTEMPLATE (0x0003)
value CDERR_REGISTERMSGFAIL (0x000C)
value CDERR_STRUCTSIZE (0x0001)
value CDM_FIRST ((WM_USER + 100))
value CDM_GETFILEPATH ((CDM_FIRST + 0x0001))
value CDM_GETFOLDERIDLIST ((CDM_FIRST + 0x0003))
value CDM_GETFOLDERPATH ((CDM_FIRST + 0x0002))
value CDM_GETSPEC ((CDM_FIRST + 0x0000))
value CDM_HIDECONTROL ((CDM_FIRST + 0x0005))
value CDM_LAST ((WM_USER + 200))
value CDM_SETCONTROLTEXT ((CDM_FIRST + 0x0004))
value CDM_SETDEFEXT ((CDM_FIRST + 0x0006))
value CDN_FILEOK ((CDN_FIRST - 0x0005))
value CDN_FIRST ((0U-601U))
value CDN_FOLDERCHANGE ((CDN_FIRST - 0x0002))
value CDN_HELP ((CDN_FIRST - 0x0004))
value CDN_INCLUDEITEM ((CDN_FIRST - 0x0007))
value CDN_INITDONE ((CDN_FIRST - 0x0000))
value CDN_LAST ((0U-699U))
value CDN_SELCHANGE ((CDN_FIRST - 0x0001))
value CDN_SHAREVIOLATION ((CDN_FIRST - 0x0003))
value CDN_TYPECHANGE ((CDN_FIRST - 0x0006))
value CDS_DISABLE_UNSAFE_MODES (0x00000200)
value CDS_ENABLE_UNSAFE_MODES (0x00000100)
value CDS_FULLSCREEN (0x00000004)
value CDS_GLOBAL (0x00000008)
value CDS_NORESET (0x10000000)
value CDS_RESET (0x40000000)
value CDS_RESET_EX (0x20000000)
value CDS_SET_PRIMARY (0x00000010)
value CDS_TEST (0x00000002)
value CDS_UPDATEREGISTRY (0x00000001)
value CDS_VIDEOPARAMETERS (0x00000020)
value CD_LBSELADD (2)
value CD_LBSELCHANGE (0)
value CD_LBSELNOITEMS (-1)
value CD_LBSELSUB (1)
value CERTSRV_E_ADMIN_DENIED_REQUEST (_HRESULT_TYPEDEF_(0x80094014L))
value CERTSRV_E_ALIGNMENT_FAULT (_HRESULT_TYPEDEF_(0x80094010L))
value CERTSRV_E_ARCHIVED_KEY_REQUIRED (_HRESULT_TYPEDEF_(0x80094804L))
value CERTSRV_E_ARCHIVED_KEY_UNEXPECTED (_HRESULT_TYPEDEF_(0x80094810L))
value CERTSRV_E_BAD_RENEWAL_CERT_ATTRIBUTE (_HRESULT_TYPEDEF_(0x8009400EL))
value CERTSRV_E_BAD_RENEWAL_SUBJECT (_HRESULT_TYPEDEF_(0x80094806L))
value CERTSRV_E_BAD_REQUESTSTATUS (_HRESULT_TYPEDEF_(0x80094003L))
value CERTSRV_E_BAD_REQUESTSUBJECT (_HRESULT_TYPEDEF_(0x80094001L))
value CERTSRV_E_BAD_REQUEST_KEY_ARCHIVAL (_HRESULT_TYPEDEF_(0x8009400CL))
value CERTSRV_E_BAD_TEMPLATE_VERSION (_HRESULT_TYPEDEF_(0x80094807L))
value CERTSRV_E_CERT_TYPE_OVERLAP (_HRESULT_TYPEDEF_(0x80094814L))
value CERTSRV_E_CORRUPT_KEY_ATTESTATION (_HRESULT_TYPEDEF_(0x8009481BL))
value CERTSRV_E_DOWNLEVEL_DC_SSL_OR_UPGRADE (_HRESULT_TYPEDEF_(0x80094013L))
value CERTSRV_E_ENCODING_LENGTH (_HRESULT_TYPEDEF_(0x80094007L))
value CERTSRV_E_ENCRYPTION_CERT_REQUIRED (_HRESULT_TYPEDEF_(0x80094018L))
value CERTSRV_E_ENROLL_DENIED (_HRESULT_TYPEDEF_(0x80094011L))
value CERTSRV_E_EXPIRED_CHALLENGE (_HRESULT_TYPEDEF_(0x8009481CL))
value CERTSRV_E_INVALID_ATTESTATION (_HRESULT_TYPEDEF_(0x80094819L))
value CERTSRV_E_INVALID_CA_CERTIFICATE (_HRESULT_TYPEDEF_(0x80094005L))
value CERTSRV_E_INVALID_EK (_HRESULT_TYPEDEF_(0x80094817L))
value CERTSRV_E_INVALID_IDBINDING (_HRESULT_TYPEDEF_(0x80094818L))
value CERTSRV_E_INVALID_REQUESTID (_HRESULT_TYPEDEF_(0x8009481EL))
value CERTSRV_E_INVALID_RESPONSE (_HRESULT_TYPEDEF_(0x8009481DL))
value CERTSRV_E_ISSUANCE_POLICY_REQUIRED (_HRESULT_TYPEDEF_(0x8009480CL))
value CERTSRV_E_KEY_ARCHIVAL_NOT_CONFIGURED (_HRESULT_TYPEDEF_(0x8009400AL))
value CERTSRV_E_KEY_ATTESTATION (_HRESULT_TYPEDEF_(0x8009481AL))
value CERTSRV_E_KEY_ATTESTATION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80094017L))
value CERTSRV_E_KEY_LENGTH (_HRESULT_TYPEDEF_(0x80094811L))
value CERTSRV_E_NO_CAADMIN_DEFINED (_HRESULT_TYPEDEF_(0x8009400DL))
value CERTSRV_E_NO_CERT_TYPE (_HRESULT_TYPEDEF_(0x80094801L))
value CERTSRV_E_NO_DB_SESSIONS (_HRESULT_TYPEDEF_(0x8009400FL))
value CERTSRV_E_NO_POLICY_SERVER (_HRESULT_TYPEDEF_(0x80094015L))
value CERTSRV_E_NO_REQUEST (_HRESULT_TYPEDEF_(0x80094002L))
value CERTSRV_E_NO_VALID_KRA (_HRESULT_TYPEDEF_(0x8009400BL))
value CERTSRV_E_PENDING_CLIENT_RESPONSE (_HRESULT_TYPEDEF_(0x80094820L))
value CERTSRV_E_PROPERTY_EMPTY (_HRESULT_TYPEDEF_(0x80094004L))
value CERTSRV_E_RENEWAL_BAD_PUBLIC_KEY (_HRESULT_TYPEDEF_(0x80094816L))
value CERTSRV_E_REQUEST_PRECERTIFICATE_MISMATCH (_HRESULT_TYPEDEF_(0x8009481FL))
value CERTSRV_E_RESTRICTEDOFFICER (_HRESULT_TYPEDEF_(0x80094009L))
value CERTSRV_E_ROLECONFLICT (_HRESULT_TYPEDEF_(0x80094008L))
value CERTSRV_E_SEC_EXT_DIRECTORY_SID_REQUIRED (_HRESULT_TYPEDEF_(0x80094821L))
value CERTSRV_E_SERVER_SUSPENDED (_HRESULT_TYPEDEF_(0x80094006L))
value CERTSRV_E_SIGNATURE_COUNT (_HRESULT_TYPEDEF_(0x8009480AL))
value CERTSRV_E_SIGNATURE_POLICY_REQUIRED (_HRESULT_TYPEDEF_(0x80094809L))
value CERTSRV_E_SIGNATURE_REJECTED (_HRESULT_TYPEDEF_(0x8009480BL))
value CERTSRV_E_SMIME_REQUIRED (_HRESULT_TYPEDEF_(0x80094805L))
value CERTSRV_E_SUBJECT_ALT_NAME_REQUIRED (_HRESULT_TYPEDEF_(0x80094803L))
value CERTSRV_E_SUBJECT_DIRECTORY_GUID_REQUIRED (_HRESULT_TYPEDEF_(0x8009480EL))
value CERTSRV_E_SUBJECT_DNS_REQUIRED (_HRESULT_TYPEDEF_(0x8009480FL))
value CERTSRV_E_SUBJECT_EMAIL_REQUIRED (_HRESULT_TYPEDEF_(0x80094812L))
value CERTSRV_E_SUBJECT_UPN_REQUIRED (_HRESULT_TYPEDEF_(0x8009480DL))
value CERTSRV_E_TEMPLATE_CONFLICT (_HRESULT_TYPEDEF_(0x80094802L))
value CERTSRV_E_TEMPLATE_DENIED (_HRESULT_TYPEDEF_(0x80094012L))
value CERTSRV_E_TEMPLATE_POLICY_REQUIRED (_HRESULT_TYPEDEF_(0x80094808L))
value CERTSRV_E_TOO_MANY_SIGNATURES (_HRESULT_TYPEDEF_(0x80094815L))
value CERTSRV_E_UNKNOWN_CERT_TYPE (_HRESULT_TYPEDEF_(0x80094813L))
value CERTSRV_E_UNSUPPORTED_CERT_TYPE (_HRESULT_TYPEDEF_(0x80094800L))
value CERTSRV_E_WEAK_SIGNATURE_OR_KEY (_HRESULT_TYPEDEF_(0x80094016L))
value CERT_ACCESS_STATE_GP_SYSTEM_STORE_FLAG (0x8)
value CERT_ACCESS_STATE_LM_SYSTEM_STORE_FLAG (0x4)
value CERT_ACCESS_STATE_PROP_ID (14)
value CERT_ACCESS_STATE_SHARED_USER_FLAG (0x10)
value CERT_ACCESS_STATE_SYSTEM_STORE_FLAG (0x2)
value CERT_ACCESS_STATE_WRITE_PERSIST_FLAG (0x1)
value CERT_AIA_URL_RETRIEVED_PROP_ID (67)
value CERT_ALT_NAME_DIRECTORY_NAME (5)
value CERT_ALT_NAME_DNS_NAME (3)
value CERT_ALT_NAME_EDI_PARTY_NAME (6)
value CERT_ALT_NAME_ENTRY_ERR_INDEX_MASK (0xFF)
value CERT_ALT_NAME_ENTRY_ERR_INDEX_SHIFT (16)
value CERT_ALT_NAME_IP_ADDRESS (8)
value CERT_ALT_NAME_OTHER_NAME (1)
value CERT_ALT_NAME_REGISTERED_ID (9)
value CERT_ALT_NAME_URL (7)
value CERT_ALT_NAME_VALUE_ERR_INDEX_MASK (0x0000FFFF)
value CERT_ALT_NAME_VALUE_ERR_INDEX_SHIFT (0)
value CERT_ARCHIVED_KEY_HASH_PROP_ID (65)
value CERT_ARCHIVED_PROP_ID (19)
value CERT_AUTHORITY_INFO_ACCESS_PROP_ID (68)
value CERT_AUTH_ROOT_AUTO_UPDATE_DISABLE_PARTIAL_CHAIN_LOGGING_FLAG (0x2)
value CERT_AUTH_ROOT_AUTO_UPDATE_DISABLE_UNTRUSTED_ROOT_LOGGING_FLAG (0x1)
value CERT_AUTH_ROOT_AUTO_UPDATE_LOCAL_MACHINE_REGPATH (CERT_AUTO_UPDATE_LOCAL_MACHINE_REGPATH)
value CERT_AUTH_ROOT_AUTO_UPDATE_ROOT_DIR_URL_VALUE_NAME (CERT_AUTO_UPDATE_ROOT_DIR_URL_VALUE_NAME)
value CERT_AUTO_ENROLL_PROP_ID (21)
value CERT_AUTO_ENROLL_RETRY_PROP_ID (66)
value CERT_AUTO_UPDATE_DISABLE_RANDOM_QUERY_STRING_FLAG (0x4)
value CERT_BACKED_UP_PROP_ID (69)
value CERT_BIOMETRIC_OID_DATA_CHOICE (2)
value CERT_BIOMETRIC_PICTURE_TYPE (0)
value CERT_BIOMETRIC_PREDEFINED_DATA_CHOICE (1)
value CERT_BIOMETRIC_SIGNATURE_TYPE (1)
value CERT_BUNDLE_CERTIFICATE (0)
value CERT_BUNDLE_CRL (1)
value CERT_CASE_INSENSITIVE_IS_RDN_ATTRS_FLAG (0x2)
value CERT_CA_DISABLE_CRL_PROP_ID (82)
value CERT_CA_OCSP_AUTHORITY_INFO_ACCESS_PROP_ID (81)
value CERT_CA_SUBJECT_FLAG (0x80)
value CERT_CEP_PROP_ID (87)
value CERT_CHAIN_AUTO_CURRENT_USER (1)
value CERT_CHAIN_AUTO_FLUSH_DISABLE_FLAG (0x00000001)
value CERT_CHAIN_AUTO_HPKP_RULE_INFO (8)
value CERT_CHAIN_AUTO_IMPERSONATED (3)
value CERT_CHAIN_AUTO_LOCAL_MACHINE (2)
value CERT_CHAIN_AUTO_LOG_CREATE_FLAG (0x00000002)
value CERT_CHAIN_AUTO_LOG_FLAGS (( CERT_CHAIN_AUTO_LOG_CREATE_FLAG | CERT_CHAIN_AUTO_LOG_FREE_FLAG | CERT_CHAIN_AUTO_LOG_FLUSH_FLAG ))
value CERT_CHAIN_AUTO_LOG_FLUSH_FLAG (0x00000008)
value CERT_CHAIN_AUTO_LOG_FREE_FLAG (0x00000004)
value CERT_CHAIN_AUTO_NETWORK_INFO (6)
value CERT_CHAIN_AUTO_PINRULE_INFO (5)
value CERT_CHAIN_AUTO_PROCESS_INFO (4)
value CERT_CHAIN_AUTO_SERIAL_LOCAL_MACHINE (7)
value CERT_CHAIN_CACHE_END_CERT (0x00000001)
value CERT_CHAIN_CACHE_ONLY_URL_RETRIEVAL (0x00000004)
value CERT_CHAIN_CRL_VALIDITY_EXT_PERIOD_HOURS_DEFAULT (12)
value CERT_CHAIN_DISABLE_AIA (0x00002000)
value CERT_CHAIN_DISABLE_ALL_EKU_WEAK_FLAG (0x00010000)
value CERT_CHAIN_DISABLE_AUTH_ROOT_AUTO_UPDATE (0x00000100)
value CERT_CHAIN_DISABLE_CODE_SIGNING_WEAK_FLAG (0x00400000)
value CERT_CHAIN_DISABLE_ECC_PARA_FLAG (0x00000010)
value CERT_CHAIN_DISABLE_FILE_HASH_WEAK_FLAG (0x00001000)
value CERT_CHAIN_DISABLE_FILE_HASH_WEAK_FLAGS (( CERT_CHAIN_DISABLE_FILE_HASH_WEAK_FLAG | CERT_CHAIN_DISABLE_MOTW_FILE_HASH_WEAK_FLAG ))
value CERT_CHAIN_DISABLE_MOTW_CODE_SIGNING_WEAK_FLAG (0x00800000)
value CERT_CHAIN_DISABLE_MOTW_FILE_HASH_WEAK_FLAG (0x00002000)
value CERT_CHAIN_DISABLE_MOTW_TIMESTAMP_HASH_WEAK_FLAG (0x00008000)
value CERT_CHAIN_DISABLE_MOTW_TIMESTAMP_WEAK_FLAG (0x08000000)
value CERT_CHAIN_DISABLE_MY_PEER_TRUST (0x00000800)
value CERT_CHAIN_DISABLE_OPT_IN_SERVER_AUTH_WEAK_FLAG (0x00040000)
value CERT_CHAIN_DISABLE_SERVER_AUTH_WEAK_FLAG (0x00100000)
value CERT_CHAIN_DISABLE_TIMESTAMP_HASH_WEAK_FLAG (0x00004000)
value CERT_CHAIN_DISABLE_TIMESTAMP_HASH_WEAK_FLAGS (( CERT_CHAIN_DISABLE_TIMESTAMP_HASH_WEAK_FLAG | CERT_CHAIN_DISABLE_MOTW_TIMESTAMP_HASH_WEAK_FLAG ))
value CERT_CHAIN_DISABLE_TIMESTAMP_WEAK_FLAG (0x04000000)
value CERT_CHAIN_DISABLE_WEAK_FLAGS (( CERT_CHAIN_DISABLE_ECC_PARA_FLAG | CERT_CHAIN_DISABLE_ALL_EKU_WEAK_FLAG | CERT_CHAIN_DISABLE_SERVER_AUTH_WEAK_FLAG | CERT_CHAIN_DISABLE_OPT_IN_SERVER_AUTH_WEAK_FLAG | CERT_CHAIN_DISABLE_CODE_SIGNING_WEAK_FLAG | CERT_CHAIN_DISABLE_MOTW_CODE_SIGNING_WEAK_FLAG | CERT_CHAIN_DISABLE_TIMESTAMP_WEAK_FLAG | CERT_CHAIN_DISABLE_MOTW_TIMESTAMP_WEAK_FLAG ))
value CERT_CHAIN_ENABLE_ALL_EKU_HYGIENE_FLAG (0x00020000)
value CERT_CHAIN_ENABLE_CACHE_AUTO_UPDATE (0x00000010)
value CERT_CHAIN_ENABLE_CODE_SIGNING_HYGIENE_FLAG (0x01000000)
value CERT_CHAIN_ENABLE_DISALLOWED_CA (0x00020000)
value CERT_CHAIN_ENABLE_HYGIENE_FLAGS (( CERT_CHAIN_ENABLE_ALL_EKU_HYGIENE_FLAG | CERT_CHAIN_ENABLE_SERVER_AUTH_HYGIENE_FLAG | CERT_CHAIN_ENABLE_CODE_SIGNING_HYGIENE_FLAG | CERT_CHAIN_ENABLE_MOTW_CODE_SIGNING_HYGIENE_FLAG | CERT_CHAIN_ENABLE_TIMESTAMP_HYGIENE_FLAG | CERT_CHAIN_ENABLE_MOTW_TIMESTAMP_HYGIENE_FLAG ))
value CERT_CHAIN_ENABLE_MOTW_CODE_SIGNING_HYGIENE_FLAG (0x02000000)
value CERT_CHAIN_ENABLE_MOTW_TIMESTAMP_HYGIENE_FLAG (0x20000000)
value CERT_CHAIN_ENABLE_ONLY_WEAK_LOGGING_FLAG (0x00000008)
value CERT_CHAIN_ENABLE_PEER_TRUST (0x00000400)
value CERT_CHAIN_ENABLE_SERVER_AUTH_HYGIENE_FLAG (0x00200000)
value CERT_CHAIN_ENABLE_SHARE_STORE (0x00000020)
value CERT_CHAIN_ENABLE_TIMESTAMP_HYGIENE_FLAG (0x10000000)
value CERT_CHAIN_ENABLE_WEAK_LOGGING_FLAG (0x00000004)
value CERT_CHAIN_ENABLE_WEAK_RSA_ROOT_FLAG (0x00000002)
value CERT_CHAIN_ENABLE_WEAK_SETTINGS_FLAG (0x80000000)
value CERT_CHAIN_EXCLUSIVE_ENABLE_CA_FLAG (0x00000001)
value CERT_CHAIN_FIND_BY_ISSUER (1)
value CERT_CHAIN_FIND_BY_ISSUER_CACHE_ONLY_FLAG (0x8000)
value CERT_CHAIN_FIND_BY_ISSUER_CACHE_ONLY_URL_FLAG (0x0004)
value CERT_CHAIN_FIND_BY_ISSUER_COMPARE_KEY_FLAG (0x0001)
value CERT_CHAIN_FIND_BY_ISSUER_COMPLEX_CHAIN_FLAG (0x0002)
value CERT_CHAIN_FIND_BY_ISSUER_LOCAL_MACHINE_FLAG (0x0008)
value CERT_CHAIN_FIND_BY_ISSUER_NO_KEY_FLAG (0x4000)
value CERT_CHAIN_HAS_MOTW (0x00004000)
value CERT_CHAIN_MAX_AIA_URL_COUNT_IN_CERT_DEFAULT (5)
value CERT_CHAIN_MAX_AIA_URL_RETRIEVAL_BYTE_COUNT_DEFAULT (100000)
value CERT_CHAIN_MAX_AIA_URL_RETRIEVAL_CERT_COUNT_DEFAULT (10)
value CERT_CHAIN_MAX_AIA_URL_RETRIEVAL_COUNT_PER_CHAIN_DEFAULT (3)
value CERT_CHAIN_MAX_SSL_TIME_UPDATED_EVENT_COUNT_DEFAULT (5)
value CERT_CHAIN_MAX_SSL_TIME_UPDATED_EVENT_COUNT_DISABLE (0xFFFFFFFF)
value CERT_CHAIN_MIN_PUB_KEY_BIT_LENGTH_DISABLE (0xFFFFFFFF)
value CERT_CHAIN_MIN_RSA_PUB_KEY_BIT_LENGTH_DEFAULT (1023)
value CERT_CHAIN_MIN_RSA_PUB_KEY_BIT_LENGTH_DISABLE (0xFFFFFFFF)
value CERT_CHAIN_MOTW_IGNORE_AFTER_TIME_WEAK_FLAG (0x40000000)
value CERT_CHAIN_MOTW_WEAK_FLAGS (( CERT_CHAIN_DISABLE_MOTW_CODE_SIGNING_WEAK_FLAG | CERT_CHAIN_DISABLE_MOTW_TIMESTAMP_WEAK_FLAG | CERT_CHAIN_ENABLE_MOTW_CODE_SIGNING_HYGIENE_FLAG | CERT_CHAIN_ENABLE_MOTW_TIMESTAMP_HYGIENE_FLAG | CERT_CHAIN_MOTW_IGNORE_AFTER_TIME_WEAK_FLAG))
value CERT_CHAIN_ONLY_ADDITIONAL_AND_AUTH_ROOT (0x00008000)
value CERT_CHAIN_OPTION_DISABLE_AIA_URL_RETRIEVAL (0x2)
value CERT_CHAIN_OPTION_ENABLE_SIA_URL_RETRIEVAL (0x4)
value CERT_CHAIN_OPT_IN_WEAK_FLAGS (( CERT_CHAIN_DISABLE_OPT_IN_SERVER_AUTH_WEAK_FLAG))
value CERT_CHAIN_OPT_IN_WEAK_SIGNATURE (0x00010000)
value CERT_CHAIN_POLICY_ALLOW_TESTROOT_FLAG (0x00008000)
value CERT_CHAIN_POLICY_ALLOW_UNKNOWN_CA_FLAG (0x00000010)
value CERT_CHAIN_POLICY_AUTHENTICODE (((LPCSTR) 2))
value CERT_CHAIN_POLICY_AUTHENTICODE_TS (((LPCSTR) 3))
value CERT_CHAIN_POLICY_BASE (((LPCSTR) 1))
value CERT_CHAIN_POLICY_BASIC_CONSTRAINTS (((LPCSTR) 5))
value CERT_CHAIN_POLICY_EV (((LPCSTR) 8))
value CERT_CHAIN_POLICY_IGNORE_ALL_NOT_TIME_VALID_FLAGS (( CERT_CHAIN_POLICY_IGNORE_NOT_TIME_VALID_FLAG | CERT_CHAIN_POLICY_IGNORE_CTL_NOT_TIME_VALID_FLAG | CERT_CHAIN_POLICY_IGNORE_NOT_TIME_NESTED_FLAG ))
value CERT_CHAIN_POLICY_IGNORE_ALL_REV_UNKNOWN_FLAGS (( CERT_CHAIN_POLICY_IGNORE_END_REV_UNKNOWN_FLAG | CERT_CHAIN_POLICY_IGNORE_CTL_SIGNER_REV_UNKNOWN_FLAG | CERT_CHAIN_POLICY_IGNORE_CA_REV_UNKNOWN_FLAG | CERT_CHAIN_POLICY_IGNORE_ROOT_REV_UNKNOWN_FLAG ))
value CERT_CHAIN_POLICY_IGNORE_CA_REV_UNKNOWN_FLAG (0x00000400)
value CERT_CHAIN_POLICY_IGNORE_CTL_NOT_TIME_VALID_FLAG (0x00000002)
value CERT_CHAIN_POLICY_IGNORE_CTL_SIGNER_REV_UNKNOWN_FLAG (0x00000200)
value CERT_CHAIN_POLICY_IGNORE_END_REV_UNKNOWN_FLAG (0x00000100)
value CERT_CHAIN_POLICY_IGNORE_INVALID_BASIC_CONSTRAINTS_FLAG (0x00000008)
value CERT_CHAIN_POLICY_IGNORE_INVALID_NAME_FLAG (0x00000040)
value CERT_CHAIN_POLICY_IGNORE_INVALID_POLICY_FLAG (0x00000080)
value CERT_CHAIN_POLICY_IGNORE_NOT_SUPPORTED_CRITICAL_EXT_FLAG (0x00002000)
value CERT_CHAIN_POLICY_IGNORE_NOT_TIME_NESTED_FLAG (0x00000004)
value CERT_CHAIN_POLICY_IGNORE_NOT_TIME_VALID_FLAG (0x00000001)
value CERT_CHAIN_POLICY_IGNORE_PEER_TRUST_FLAG (0x00001000)
value CERT_CHAIN_POLICY_IGNORE_ROOT_REV_UNKNOWN_FLAG (0x00000800)
value CERT_CHAIN_POLICY_IGNORE_WEAK_SIGNATURE_FLAG (0x08000000)
value CERT_CHAIN_POLICY_IGNORE_WRONG_USAGE_FLAG (0x00000020)
value CERT_CHAIN_POLICY_MICROSOFT_ROOT (((LPCSTR) 7))
value CERT_CHAIN_POLICY_NT_AUTH (((LPCSTR) 6))
value CERT_CHAIN_POLICY_SSL (((LPCSTR) 4))
value CERT_CHAIN_POLICY_SSL_HPKP_HEADER (((LPCSTR) 10))
value CERT_CHAIN_POLICY_SSL_KEY_PIN (((LPCSTR) 12))
value CERT_CHAIN_POLICY_SSL_KEY_PIN_MISMATCH_ERROR (-2)
value CERT_CHAIN_POLICY_SSL_KEY_PIN_MISMATCH_WARNING (2)
value CERT_CHAIN_POLICY_SSL_KEY_PIN_MITM_ERROR (-1)
value CERT_CHAIN_POLICY_SSL_KEY_PIN_MITM_WARNING (1)
value CERT_CHAIN_POLICY_SSL_KEY_PIN_SUCCESS (0)
value CERT_CHAIN_POLICY_THIRD_PARTY_ROOT (((LPCSTR) 11))
value CERT_CHAIN_POLICY_TRUST_TESTROOT_FLAG (0x00004000)
value CERT_CHAIN_RETURN_LOWER_QUALITY_CONTEXTS (0x00000080)
value CERT_CHAIN_REVOCATION_ACCUMULATIVE_TIMEOUT (0x08000000)
value CERT_CHAIN_REVOCATION_CHECK_CACHE_ONLY (0x80000000)
value CERT_CHAIN_REVOCATION_CHECK_CHAIN (0x20000000)
value CERT_CHAIN_REVOCATION_CHECK_CHAIN_EXCLUDE_ROOT (0x40000000)
value CERT_CHAIN_REVOCATION_CHECK_END_CERT (0x10000000)
value CERT_CHAIN_REVOCATION_CHECK_OCSP_CERT (0x04000000)
value CERT_CHAIN_STRONG_SIGN_DISABLE_END_CHECK_FLAG (0x00000001)
value CERT_CHAIN_THREAD_STORE_SYNC (0x00000002)
value CERT_CHAIN_TIMESTAMP_TIME (0x00000200)
value CERT_CHAIN_USE_LOCAL_MACHINE_STORE (0x00000008)
value CERT_CLOSE_STORE_CHECK_FLAG (0x00000002)
value CERT_CLOSE_STORE_FORCE_FLAG (0x00000001)
value CERT_CLR_DELETE_KEY_PROP_ID (125)
value CERT_COMPARE_ANY (0)
value CERT_COMPARE_ATTR (3)
value CERT_COMPARE_CERT_ID (16)
value CERT_COMPARE_CROSS_CERT_DIST_POINTS (17)
value CERT_COMPARE_CTL_USAGE (CERT_COMPARE_ENHKEY_USAGE)
value CERT_COMPARE_ENHKEY_USAGE (10)
value CERT_COMPARE_EXISTING (13)
value CERT_COMPARE_HASH (CERT_COMPARE_SHA1_HASH)
value CERT_COMPARE_HASH_STR (20)
value CERT_COMPARE_HAS_PRIVATE_KEY (21)
value CERT_COMPARE_ISSUER_OF (12)
value CERT_COMPARE_KEY_IDENTIFIER (15)
value CERT_COMPARE_KEY_SPEC (9)
value CERT_COMPARE_MASK (0xFFFF)
value CERT_COMPARE_NAME (2)
value CERT_COMPARE_NAME_STR_A (7)
value CERT_COMPARE_NAME_STR_W (8)
value CERT_COMPARE_PROPERTY (5)
value CERT_COMPARE_PUBLIC_KEY (6)
value CERT_COMPARE_SHIFT (16)
value CERT_COMPARE_SIGNATURE_HASH (14)
value CERT_COMPARE_SUBJECT_CERT (11)
value CERT_COMPARE_SUBJECT_INFO_ACCESS (19)
value CERT_CONTEXT_REVOCATION_TYPE (1)
value CERT_CREATE_CONTEXT_NOCOPY_FLAG (0x1)
value CERT_CREATE_CONTEXT_NO_ENTRY_FLAG (0x8)
value CERT_CREATE_CONTEXT_NO_HCRYPTMSG_FLAG (0x4)
value CERT_CREATE_CONTEXT_SORTED_FLAG (0x2)
value CERT_CREATE_SELFSIGN_NO_KEY_INFO (2)
value CERT_CREATE_SELFSIGN_NO_SIGN (1)
value CERT_CRL_SIGN_KEY_USAGE (0x02)
value CERT_CROSS_CERT_DIST_POINTS_PROP_ID (23)
value CERT_CTL_USAGE_PROP_ID (CERT_ENHKEY_USAGE_PROP_ID)
value CERT_DATA_ENCIPHERMENT_KEY_USAGE (0x10)
value CERT_DATE_STAMP_PROP_ID (27)
value CERT_DECIPHER_ONLY_KEY_USAGE (0x80)
value CERT_DESCRIPTION_PROP_ID (13)
value CERT_DIGITAL_SIGNATURE_KEY_USAGE (0x80)
value CERT_DISALLOWED_CA_FILETIME_PROP_ID (128)
value CERT_DISALLOWED_ENHKEY_USAGE_PROP_ID (122)
value CERT_DISALLOWED_FILETIME_PROP_ID (104)
value CERT_DSS_R_LEN (20)
value CERT_DSS_SIGNATURE_LEN ((CERT_DSS_R_LEN + CERT_DSS_S_LEN))
value CERT_DSS_S_LEN (20)
value CERT_EFS_PROP_ID (17)
value CERT_ENCIPHER_ONLY_KEY_USAGE (0x01)
value CERT_ENCODING_TYPE_MASK (0x0000FFFF)
value CERT_END_ENTITY_SUBJECT_FLAG (0x40)
value CERT_ENHKEY_USAGE_PROP_ID (9)
value CERT_ENROLLMENT_PROP_ID (26)
value CERT_EXCLUDED_SUBTREE_BIT (0x80000000L)
value CERT_EXTENDED_ERROR_INFO_PROP_ID (30)
value CERT_E_CHAINING (_HRESULT_TYPEDEF_(0x800B010AL))
value CERT_E_CN_NO_MATCH (_HRESULT_TYPEDEF_(0x800B010FL))
value CERT_E_CRITICAL (_HRESULT_TYPEDEF_(0x800B0105L))
value CERT_E_EXPIRED (_HRESULT_TYPEDEF_(0x800B0101L))
value CERT_E_INVALID_NAME (_HRESULT_TYPEDEF_(0x800B0114L))
value CERT_E_INVALID_POLICY (_HRESULT_TYPEDEF_(0x800B0113L))
value CERT_E_ISSUERCHAINING (_HRESULT_TYPEDEF_(0x800B0107L))
value CERT_E_MALFORMED (_HRESULT_TYPEDEF_(0x800B0108L))
value CERT_E_PATHLENCONST (_HRESULT_TYPEDEF_(0x800B0104L))
value CERT_E_PURPOSE (_HRESULT_TYPEDEF_(0x800B0106L))
value CERT_E_REVOCATION_FAILURE (_HRESULT_TYPEDEF_(0x800B010EL))
value CERT_E_REVOKED (_HRESULT_TYPEDEF_(0x800B010CL))
value CERT_E_ROLE (_HRESULT_TYPEDEF_(0x800B0103L))
value CERT_E_UNTRUSTEDCA (_HRESULT_TYPEDEF_(0x800B0112L))
value CERT_E_UNTRUSTEDROOT (_HRESULT_TYPEDEF_(0x800B0109L))
value CERT_E_UNTRUSTEDTESTROOT (_HRESULT_TYPEDEF_(0x800B010DL))
value CERT_E_VALIDITYPERIODNESTING (_HRESULT_TYPEDEF_(0x800B0102L))
value CERT_E_WRONG_USAGE (_HRESULT_TYPEDEF_(0x800B0110L))
value CERT_FILE_HASH_USE_TYPE (1)
value CERT_FILE_STORE_COMMIT_ENABLE_FLAG (0x10000)
value CERT_FIND_CTL_USAGE (CERT_FIND_ENHKEY_USAGE)
value CERT_FIND_EXT_ONLY_CTL_USAGE_FLAG (CERT_FIND_EXT_ONLY_ENHKEY_USAGE_FLAG)
value CERT_FIND_EXT_ONLY_ENHKEY_USAGE_FLAG (0x2)
value CERT_FIND_HASH (CERT_FIND_SHA1_HASH)
value CERT_FIND_ISSUER_STR (CERT_FIND_ISSUER_STR_W)
value CERT_FIND_NO_CTL_USAGE_FLAG (CERT_FIND_NO_ENHKEY_USAGE_FLAG)
value CERT_FIND_NO_ENHKEY_USAGE_FLAG (0x8)
value CERT_FIND_OPTIONAL_CTL_USAGE_FLAG (CERT_FIND_OPTIONAL_ENHKEY_USAGE_FLAG)
value CERT_FIND_OPTIONAL_ENHKEY_USAGE_FLAG (0x1)
value CERT_FIND_OR_CTL_USAGE_FLAG (CERT_FIND_OR_ENHKEY_USAGE_FLAG)
value CERT_FIND_OR_ENHKEY_USAGE_FLAG (0x10)
value CERT_FIND_PROP_ONLY_CTL_USAGE_FLAG (CERT_FIND_PROP_ONLY_ENHKEY_USAGE_FLAG)
value CERT_FIND_PROP_ONLY_ENHKEY_USAGE_FLAG (0x4)
value CERT_FIND_SUBJECT_STR (CERT_FIND_SUBJECT_STR_W)
value CERT_FIND_VALID_CTL_USAGE_FLAG (CERT_FIND_VALID_ENHKEY_USAGE_FLAG)
value CERT_FIND_VALID_ENHKEY_USAGE_FLAG (0x20)
value CERT_FIRST_RESERVED_PROP_ID (129)
value CERT_FIRST_USER_PROP_ID (0x00008000)
value CERT_FORTEZZA_DATA_PROP_ID (18)
value CERT_FRIENDLY_NAME_PROP_ID (11)
value CERT_HASH_PROP_ID (CERT_SHA1_HASH_PROP_ID)
value CERT_HCRYPTPROV_OR_NCRYPT_KEY_HANDLE_PROP_ID (79)
value CERT_HCRYPTPROV_TRANSFER_PROP_ID (100)
value CERT_ID_ISSUER_SERIAL_NUMBER (1)
value CERT_ID_KEY_IDENTIFIER (2)
value CERT_INFO_EXTENSION_FLAG (11)
value CERT_INFO_ISSUER_FLAG (4)
value CERT_INFO_ISSUER_UNIQUE_ID_FLAG (9)
value CERT_INFO_NOT_AFTER_FLAG (6)
value CERT_INFO_NOT_BEFORE_FLAG (5)
value CERT_INFO_SERIAL_NUMBER_FLAG (2)
value CERT_INFO_SIGNATURE_ALGORITHM_FLAG (3)
value CERT_INFO_SUBJECT_FLAG (7)
value CERT_INFO_SUBJECT_PUBLIC_KEY_INFO_FLAG (8)
value CERT_INFO_SUBJECT_UNIQUE_ID_FLAG (10)
value CERT_INFO_VERSION_FLAG (1)
value CERT_ISOLATED_KEY_PROP_ID (118)
value CERT_ISSUER_CHAIN_PUB_KEY_CNG_ALG_BIT_LENGTH_PROP_ID (96)
value CERT_ISSUER_CHAIN_SIGN_HASH_CNG_ALG_PROP_ID (95)
value CERT_ISSUER_PUB_KEY_BIT_LENGTH_PROP_ID (94)
value CERT_KEY_AGREEMENT_KEY_USAGE (0x08)
value CERT_KEY_CERT_SIGN_KEY_USAGE (0x04)
value CERT_KEY_CLASSIFICATION_PROP_ID (120)
value CERT_KEY_CONTEXT_PROP_ID (5)
value CERT_KEY_ENCIPHERMENT_KEY_USAGE (0x20)
value CERT_KEY_IDENTIFIER_PROP_ID (20)
value CERT_KEY_PROV_HANDLE_PROP_ID (1)
value CERT_KEY_PROV_INFO_PROP_ID (2)
value CERT_KEY_REPAIR_ATTEMPTED_PROP_ID (103)
value CERT_KEY_SPEC_PROP_ID (6)
value CERT_LAST_RESERVED_PROP_ID (0x00007FFF)
value CERT_LAST_USER_PROP_ID (0x0000FFFF)
value CERT_LDAP_STORE_AREC_EXCLUSIVE_FLAG (0x20000)
value CERT_LDAP_STORE_OPENED_FLAG (0x40000)
value CERT_LDAP_STORE_SIGN_FLAG (0x10000)
value CERT_LDAP_STORE_UNBIND_FLAG (0x80000)
value CERT_LOGOTYPE_BITS_IMAGE_RESOLUTION_CHOICE (1)
value CERT_LOGOTYPE_COLOR_IMAGE_INFO_CHOICE (2)
value CERT_LOGOTYPE_DIRECT_INFO_CHOICE (1)
value CERT_LOGOTYPE_GRAY_SCALE_IMAGE_INFO_CHOICE (1)
value CERT_LOGOTYPE_INDIRECT_INFO_CHOICE (2)
value CERT_LOGOTYPE_NO_IMAGE_RESOLUTION_CHOICE (0)
value CERT_LOGOTYPE_TABLE_SIZE_IMAGE_RESOLUTION_CHOICE (2)
value CERT_NAME_ATTR_TYPE (3)
value CERT_NAME_DNS_TYPE (6)
value CERT_NAME_EMAIL_TYPE (1)
value CERT_NAME_FRIENDLY_DISPLAY_TYPE (5)
value CERT_NAME_ISSUER_FLAG (0x1)
value CERT_NAME_RDN_TYPE (2)
value CERT_NAME_SEARCH_ALL_NAMES_FLAG (0x2)
value CERT_NAME_SIMPLE_DISPLAY_TYPE (4)
value CERT_NAME_STR_COMMA_FLAG (0x04000000)
value CERT_NAME_STR_CRLF_FLAG (0x08000000)
value CERT_NAME_STR_ENABLE_PUNYCODE_FLAG (0x00200000)
value CERT_NAME_STR_FORWARD_FLAG (0x01000000)
value CERT_NAME_STR_NO_PLUS_FLAG (0x20000000)
value CERT_NAME_STR_NO_QUOTING_FLAG (0x10000000)
value CERT_NAME_STR_REVERSE_FLAG (0x02000000)
value CERT_NAME_STR_SEMICOLON_FLAG (0x40000000)
value CERT_NAME_UPN_TYPE (8)
value CERT_NAME_URL_TYPE (7)
value CERT_NCRYPT_KEY_HANDLE_PROP_ID (78)
value CERT_NCRYPT_KEY_HANDLE_TRANSFER_PROP_ID (99)
value CERT_NCRYPT_KEY_SPEC (0xFFFFFFFF)
value CERT_NEW_KEY_PROP_ID (74)
value CERT_NEXT_UPDATE_LOCATION_PROP_ID (10)
value CERT_NONCOMPLIANT_ROOT_URL_PROP_ID (123)
value CERT_NON_REPUDIATION_KEY_USAGE (0x40)
value CERT_NOT_BEFORE_ENHKEY_USAGE_PROP_ID (127)
value CERT_NOT_BEFORE_FILETIME_PROP_ID (126)
value CERT_NO_AUTO_EXPIRE_CHECK_PROP_ID (77)
value CERT_NO_EXPIRE_NOTIFICATION_PROP_ID (97)
value CERT_OCSP_CACHE_PREFIX_PROP_ID (75)
value CERT_OCSP_MUST_STAPLE_PROP_ID (121)
value CERT_OCSP_RESPONSE_PROP_ID (70)
value CERT_OFFLINE_CRL_SIGN_KEY_USAGE (0x02)
value CERT_OID_NAME_STR (2)
value CERT_PHYSICAL_STORE_ADD_ENABLE_FLAG (0x1)
value CERT_PHYSICAL_STORE_INSERT_COMPUTER_NAME_ENABLE_FLAG (0x8)
value CERT_PHYSICAL_STORE_OPEN_DISABLE_FLAG (0x2)
value CERT_PHYSICAL_STORE_PREDEFINED_ENUM_FLAG (0x1)
value CERT_PHYSICAL_STORE_REMOTE_OPEN_DISABLE_FLAG (0x4)
value CERT_PROT_ROOT_DISABLE_CURRENT_USER_FLAG (0x1)
value CERT_PROT_ROOT_DISABLE_LM_AUTH_FLAG (0x8)
value CERT_PROT_ROOT_DISABLE_NOT_DEFINED_NAME_CONSTRAINT_FLAG (0x20)
value CERT_PROT_ROOT_DISABLE_NT_AUTH_REQUIRED_FLAG (0x10)
value CERT_PROT_ROOT_DISABLE_PEER_TRUST (0x10000)
value CERT_PROT_ROOT_INHIBIT_ADD_AT_INIT_FLAG (0x2)
value CERT_PROT_ROOT_INHIBIT_PURGE_LM_FLAG (0x4)
value CERT_PROT_ROOT_ONLY_LM_GPT_FLAG (0x8)
value CERT_PUBKEY_ALG_PARA_PROP_ID (22)
value CERT_PUBKEY_HASH_RESERVED_PROP_ID (8)
value CERT_PUB_KEY_CNG_ALG_BIT_LENGTH_PROP_ID (93)
value CERT_PVK_FILE_PROP_ID (12)
value CERT_QUERY_CONTENT_CERT (1)
value CERT_QUERY_CONTENT_CERT_PAIR (13)
value CERT_QUERY_CONTENT_CRL (3)
value CERT_QUERY_CONTENT_CTL (2)
value CERT_QUERY_CONTENT_FLAG_ALL (( CERT_QUERY_CONTENT_FLAG_CERT | CERT_QUERY_CONTENT_FLAG_CTL | CERT_QUERY_CONTENT_FLAG_CRL | CERT_QUERY_CONTENT_FLAG_SERIALIZED_STORE | CERT_QUERY_CONTENT_FLAG_SERIALIZED_CERT | CERT_QUERY_CONTENT_FLAG_SERIALIZED_CTL | CERT_QUERY_CONTENT_FLAG_SERIALIZED_CRL | CERT_QUERY_CONTENT_FLAG_PKCS7_SIGNED | CERT_QUERY_CONTENT_FLAG_PKCS7_UNSIGNED | CERT_QUERY_CONTENT_FLAG_PKCS7_SIGNED_EMBED | CERT_QUERY_CONTENT_FLAG_PKCS10 | CERT_QUERY_CONTENT_FLAG_PFX | CERT_QUERY_CONTENT_FLAG_CERT_PAIR ))
value CERT_QUERY_CONTENT_FLAG_ALL_ISSUER_CERT (( CERT_QUERY_CONTENT_FLAG_CERT | CERT_QUERY_CONTENT_FLAG_SERIALIZED_STORE | CERT_QUERY_CONTENT_FLAG_SERIALIZED_CERT | CERT_QUERY_CONTENT_FLAG_PKCS7_SIGNED | CERT_QUERY_CONTENT_FLAG_PKCS7_UNSIGNED ))
value CERT_QUERY_CONTENT_PFX (12)
value CERT_QUERY_CONTENT_PFX_AND_LOAD (14)
value CERT_QUERY_CONTENT_SERIALIZED_CERT (5)
value CERT_QUERY_CONTENT_SERIALIZED_CRL (7)
value CERT_QUERY_CONTENT_SERIALIZED_CTL (6)
value CERT_QUERY_CONTENT_SERIALIZED_STORE (4)
value CERT_QUERY_FORMAT_ASN_ASCII_HEX_ENCODED (3)
value CERT_QUERY_FORMAT_BINARY (1)
value CERT_QUERY_FORMAT_FLAG_ALL (( CERT_QUERY_FORMAT_FLAG_BINARY | CERT_QUERY_FORMAT_FLAG_BASE64_ENCODED | CERT_QUERY_FORMAT_FLAG_ASN_ASCII_HEX_ENCODED ))
value CERT_QUERY_OBJECT_BLOB (0x00000002)
value CERT_QUERY_OBJECT_FILE (0x00000001)
value CERT_RDN_ANY_TYPE (0)
value CERT_RDN_BMP_STRING (12)
value CERT_RDN_DISABLE_CHECK_TYPE_FLAG (0x40000000)
value CERT_RDN_ENABLE_PUNYCODE_FLAG (0x02000000)
value CERT_RDN_ENCODED_BLOB (1)
value CERT_RDN_FLAGS_MASK (0xFF000000)
value CERT_RDN_GENERAL_STRING (10)
value CERT_RDN_GRAPHIC_STRING (8)
value CERT_RDN_NUMERIC_STRING (3)
value CERT_RDN_OCTET_STRING (2)
value CERT_RDN_PRINTABLE_STRING (4)
value CERT_RDN_TELETEX_STRING (5)
value CERT_RDN_TYPE_MASK (0x000000FF)
value CERT_RDN_UNICODE_STRING (12)
value CERT_RDN_UNIVERSAL_STRING (11)
value CERT_RDN_VIDEOTEX_STRING (6)
value CERT_RDN_VISIBLE_STRING (9)
value CERT_REGISTRY_STORE_CLIENT_GPT_FLAG (0x80000000)
value CERT_REGISTRY_STORE_EXTERNAL_FLAG (0x100000)
value CERT_REGISTRY_STORE_LM_GPT_FLAG (0x01000000)
value CERT_REGISTRY_STORE_MY_IE_DIRTY_FLAG (0x80000)
value CERT_REGISTRY_STORE_REMOTE_FLAG (0x10000)
value CERT_REGISTRY_STORE_ROAMING_FLAG (0x40000)
value CERT_REGISTRY_STORE_SERIALIZED_FLAG (0x20000)
value CERT_RENEWAL_PROP_ID (64)
value CERT_REQUEST_ORIGINATOR_PROP_ID (71)
value CERT_RETRIEVE_BIOMETRIC_PICTURE_TYPE ((CERT_RETRIEVE_BIOMETRIC_PREDEFINED_BASE_TYPE + CERT_BIOMETRIC_PICTURE_TYPE))
value CERT_RETRIEVE_BIOMETRIC_PREDEFINED_BASE_TYPE (((LPCSTR) 1000))
value CERT_RETRIEVE_BIOMETRIC_SIGNATURE_TYPE ((CERT_RETRIEVE_BIOMETRIC_PREDEFINED_BASE_TYPE + CERT_BIOMETRIC_SIGNATURE_TYPE))
value CERT_RETRIEVE_COMMUNITY_LOGO (((LPCSTR) 3))
value CERT_RETRIEVE_ISSUER_LOGO (((LPCSTR) 1))
value CERT_RETRIEVE_SUBJECT_LOGO (((LPCSTR) 2))
value CERT_ROOT_PROGRAM_CERT_POLICIES_PROP_ID (83)
value CERT_ROOT_PROGRAM_CHAIN_POLICIES_PROP_ID (105)
value CERT_ROOT_PROGRAM_FLAG_ADDRESS (0x08)
value CERT_ROOT_PROGRAM_FLAG_LSC (0x40)
value CERT_ROOT_PROGRAM_FLAG_ORG (0x80)
value CERT_ROOT_PROGRAM_FLAG_OU (0x10)
value CERT_ROOT_PROGRAM_FLAG_SUBJECT_LOGO (0x20)
value CERT_ROOT_PROGRAM_NAME_CONSTRAINTS_PROP_ID (84)
value CERT_SCARD_PIN_ID_PROP_ID (90)
value CERT_SCARD_PIN_INFO_PROP_ID (91)
value CERT_SCEP_CA_CERT_PROP_ID (111)
value CERT_SCEP_ENCRYPT_HASH_CNG_ALG_PROP_ID (114)
value CERT_SCEP_FLAGS_PROP_ID (115)
value CERT_SCEP_GUID_PROP_ID (116)
value CERT_SCEP_NONCE_PROP_ID (113)
value CERT_SCEP_RA_ENCRYPTION_CERT_PROP_ID (110)
value CERT_SCEP_RA_SIGNATURE_CERT_PROP_ID (109)
value CERT_SCEP_SERVER_CERTS_PROP_ID (108)
value CERT_SCEP_SIGNER_CERT_PROP_ID (112)
value CERT_SELECT_ALLOW_DUPLICATES (0x00000080)
value CERT_SELECT_ALLOW_EXPIRED (0x00000001)
value CERT_SELECT_BY_ENHKEY_USAGE (1)
value CERT_SELECT_BY_EXTENSION (5)
value CERT_SELECT_BY_FRIENDLYNAME (13)
value CERT_SELECT_BY_ISSUER_ATTR (7)
value CERT_SELECT_BY_ISSUER_DISPLAYNAME (12)
value CERT_SELECT_BY_ISSUER_NAME (9)
value CERT_SELECT_BY_KEY_USAGE (2)
value CERT_SELECT_BY_POLICY_OID (3)
value CERT_SELECT_BY_PROV_NAME (4)
value CERT_SELECT_BY_PUBLIC_KEY (10)
value CERT_SELECT_BY_SUBJECT_ATTR (8)
value CERT_SELECT_BY_SUBJECT_HOST_NAME (6)
value CERT_SELECT_BY_THUMBPRINT (14)
value CERT_SELECT_BY_TLS_SIGNATURES (11)
value CERT_SELECT_DISALLOW_SELFSIGNED (0x00000004)
value CERT_SELECT_HARDWARE_ONLY (0x00000040)
value CERT_SELECT_HAS_KEY_FOR_KEY_EXCHANGE (0x00000020)
value CERT_SELECT_HAS_KEY_FOR_SIGNATURE (0x00000010)
value CERT_SELECT_HAS_PRIVATE_KEY (0x00000008)
value CERT_SELECT_IGNORE_AUTOSELECT (0x00000100)
value CERT_SELECT_LAST (CERT_SELECT_BY_TLS_SIGNATURES)
value CERT_SELECT_MAX_PARA (500)
value CERT_SELECT_TRUSTED_ROOT (0x00000002)
value CERT_SEND_AS_TRUSTED_ISSUER_PROP_ID (102)
value CERT_SERIALIZABLE_KEY_CONTEXT_PROP_ID (117)
value CERT_SERIAL_CHAIN_PROP_ID (119)
value CERT_SERVER_OCSP_RESPONSE_ASYNC_FLAG (0x00000001)
value CERT_SERVER_OCSP_RESPONSE_OPEN_PARA_READ_FLAG (0x00000001)
value CERT_SERVER_OCSP_RESPONSE_OPEN_PARA_WRITE_FLAG (0x00000002)
value CERT_SET_KEY_CONTEXT_PROP_ID (0x00000001)
value CERT_SET_KEY_PROV_HANDLE_PROP_ID (0x00000001)
value CERT_SET_PROPERTY_IGNORE_PERSIST_ERROR_FLAG (0x80000000)
value CERT_SET_PROPERTY_INHIBIT_PERSIST_FLAG (0x40000000)
value CERT_SIGNATURE_HASH_PROP_ID (15)
value CERT_SIGN_HASH_CNG_ALG_PROP_ID (89)
value CERT_SIMPLE_NAME_STR (1)
value CERT_SMART_CARD_DATA_PROP_ID (16)
value CERT_SMART_CARD_READER_NON_REMOVABLE_PROP_ID (106)
value CERT_SMART_CARD_READER_PROP_ID (101)
value CERT_SMART_CARD_ROOT_INFO_PROP_ID (76)
value CERT_SOURCE_LOCATION_PROP_ID (72)
value CERT_SOURCE_URL_PROP_ID (73)
value CERT_SRV_OCSP_RESP_MIN_SYNC_CERT_FILE_SECONDS_DEFAULT (5)
value CERT_STORE_ADD_ALWAYS (4)
value CERT_STORE_ADD_NEW (1)
value CERT_STORE_ADD_NEWER (6)
value CERT_STORE_ADD_NEWER_INHERIT_PROPERTIES (7)
value CERT_STORE_ADD_REPLACE_EXISTING (3)
value CERT_STORE_ADD_REPLACE_EXISTING_INHERIT_PROPERTIES (5)
value CERT_STORE_ADD_USE_EXISTING (2)
value CERT_STORE_BACKUP_RESTORE_FLAG (0x00000800)
value CERT_STORE_BASE_CRL_FLAG (0x00000100)
value CERT_STORE_CERTIFICATE_CONTEXT (1)
value CERT_STORE_CREATE_NEW_FLAG (0x00002000)
value CERT_STORE_CRL_CONTEXT (2)
value CERT_STORE_CTL_CONTEXT (3)
value CERT_STORE_CTRL_AUTO_RESYNC (4)
value CERT_STORE_CTRL_CANCEL_NOTIFY (5)
value CERT_STORE_CTRL_COMMIT (3)
value CERT_STORE_CTRL_COMMIT_CLEAR_FLAG (0x2)
value CERT_STORE_CTRL_COMMIT_FORCE_FLAG (0x1)
value CERT_STORE_CTRL_INHIBIT_DUPLICATE_HANDLE_FLAG (0x1)
value CERT_STORE_CTRL_NOTIFY_CHANGE (2)
value CERT_STORE_CTRL_RESYNC (1)
value CERT_STORE_DEFER_CLOSE_UNTIL_LAST_FREE_FLAG (0x00000004)
value CERT_STORE_DELETE_FLAG (0x00000010)
value CERT_STORE_DELTA_CRL_FLAG (0x00000200)
value CERT_STORE_ENUM_ARCHIVED_FLAG (0x00000200)
value CERT_STORE_LOCALIZED_NAME_PROP_ID (0x1000)
value CERT_STORE_MANIFOLD_FLAG (0x00000100)
value CERT_STORE_MAXIMUM_ALLOWED_FLAG (0x00001000)
value CERT_STORE_NO_CRL_FLAG (0x00010000)
value CERT_STORE_NO_CRYPT_RELEASE_FLAG (0x00000001)
value CERT_STORE_NO_ISSUER_FLAG (0x00020000)
value CERT_STORE_OPEN_EXISTING_FLAG (0x00004000)
value CERT_STORE_PROV_CLOSE_FUNC (0)
value CERT_STORE_PROV_COLLECTION (((LPCSTR) 11))
value CERT_STORE_PROV_CONTROL_FUNC (13)
value CERT_STORE_PROV_DELETED_FLAG (0x2)
value CERT_STORE_PROV_DELETE_CERT_FUNC (3)
value CERT_STORE_PROV_DELETE_CRL_FUNC (7)
value CERT_STORE_PROV_DELETE_CTL_FUNC (11)
value CERT_STORE_PROV_EXTERNAL_FLAG (0x1)
value CERT_STORE_PROV_FILE (((LPCSTR) 3))
value CERT_STORE_PROV_FILENAME (CERT_STORE_PROV_FILENAME_W)
value CERT_STORE_PROV_FILENAME_A (((LPCSTR) 7))
value CERT_STORE_PROV_FILENAME_W (((LPCSTR) 8))
value CERT_STORE_PROV_FIND_CERT_FUNC (14)
value CERT_STORE_PROV_FIND_CRL_FUNC (17)
value CERT_STORE_PROV_FIND_CTL_FUNC (20)
value CERT_STORE_PROV_FREE_FIND_CERT_FUNC (15)
value CERT_STORE_PROV_FREE_FIND_CRL_FUNC (18)
value CERT_STORE_PROV_FREE_FIND_CTL_FUNC (21)
value CERT_STORE_PROV_GET_CERT_PROPERTY_FUNC (16)
value CERT_STORE_PROV_GET_CRL_PROPERTY_FUNC (19)
value CERT_STORE_PROV_GET_CTL_PROPERTY_FUNC (22)
value CERT_STORE_PROV_GP_SYSTEM_STORE_FLAG (0x20)
value CERT_STORE_PROV_LDAP (CERT_STORE_PROV_LDAP_W)
value CERT_STORE_PROV_LDAP_W (((LPCSTR) 16))
value CERT_STORE_PROV_LM_SYSTEM_STORE_FLAG (0x10)
value CERT_STORE_PROV_MEMORY (((LPCSTR) 2))
value CERT_STORE_PROV_MSG (((LPCSTR) 1))
value CERT_STORE_PROV_NO_PERSIST_FLAG (0x4)
value CERT_STORE_PROV_PHYSICAL (CERT_STORE_PROV_PHYSICAL_W)
value CERT_STORE_PROV_PHYSICAL_W (((LPCSTR) 14))
value CERT_STORE_PROV_READ_CERT_FUNC (1)
value CERT_STORE_PROV_READ_CRL_FUNC (5)
value CERT_STORE_PROV_READ_CTL_FUNC (9)
value CERT_STORE_PROV_REG (((LPCSTR) 4))
value CERT_STORE_PROV_SERIALIZED (((LPCSTR) 6))
value CERT_STORE_PROV_SET_CERT_PROPERTY_FUNC (4)
value CERT_STORE_PROV_SET_CRL_PROPERTY_FUNC (8)
value CERT_STORE_PROV_SET_CTL_PROPERTY_FUNC (12)
value CERT_STORE_PROV_SHARED_USER_FLAG (0x40)
value CERT_STORE_PROV_SMART_CARD (CERT_STORE_PROV_SMART_CARD_W)
value CERT_STORE_PROV_SMART_CARD_W (((LPCSTR) 15))
value CERT_STORE_PROV_SYSTEM (CERT_STORE_PROV_SYSTEM_W)
value CERT_STORE_PROV_SYSTEM_A (((LPCSTR) 9))
value CERT_STORE_PROV_SYSTEM_REGISTRY (CERT_STORE_PROV_SYSTEM_REGISTRY_W)
value CERT_STORE_PROV_SYSTEM_REGISTRY_A (((LPCSTR) 12))
value CERT_STORE_PROV_SYSTEM_REGISTRY_W (((LPCSTR) 13))
value CERT_STORE_PROV_SYSTEM_STORE_FLAG (0x8)
value CERT_STORE_PROV_SYSTEM_W (((LPCSTR) 10))
value CERT_STORE_PROV_WRITE_ADD_FLAG (0x1)
value CERT_STORE_PROV_WRITE_CERT_FUNC (2)
value CERT_STORE_PROV_WRITE_CRL_FUNC (6)
value CERT_STORE_PROV_WRITE_CTL_FUNC (10)
value CERT_STORE_READONLY_FLAG (0x00008000)
value CERT_STORE_REVOCATION_FLAG (0x00000004)
value CERT_STORE_SAVE_AS_STORE (1)
value CERT_STORE_SAVE_TO_FILE (1)
value CERT_STORE_SAVE_TO_FILENAME (CERT_STORE_SAVE_TO_FILENAME_W)
value CERT_STORE_SAVE_TO_FILENAME_A (3)
value CERT_STORE_SAVE_TO_FILENAME_W (4)
value CERT_STORE_SAVE_TO_MEMORY (2)
value CERT_STORE_SET_LOCALIZED_NAME_FLAG (0x00000002)
value CERT_STORE_SHARE_CONTEXT_FLAG (0x00000080)
value CERT_STORE_SHARE_STORE_FLAG (0x00000040)
value CERT_STORE_SIGNATURE_FLAG (0x00000001)
value CERT_STORE_TIME_VALIDITY_FLAG (0x00000002)
value CERT_STORE_UNSAFE_PHYSICAL_FLAG (0x00000020)
value CERT_STORE_UPDATE_KEYID_FLAG (0x00000400)
value CERT_STRONG_SIGN_ENABLE_CRL_CHECK (0x1)
value CERT_STRONG_SIGN_ENABLE_OCSP_CHECK (0x2)
value CERT_STRONG_SIGN_OID_INFO_CHOICE (2)
value CERT_STRONG_SIGN_SERIALIZED_INFO_CHOICE (1)
value CERT_SUBJECT_DISABLE_CRL_PROP_ID (86)
value CERT_SUBJECT_INFO_ACCESS_PROP_ID (80)
value CERT_SUBJECT_OCSP_AUTHORITY_INFO_ACCESS_PROP_ID (85)
value CERT_SUBJECT_PUB_KEY_BIT_LENGTH_PROP_ID (92)
value CERT_SYSTEM_STORE_CURRENT_SERVICE_ID (4)
value CERT_SYSTEM_STORE_CURRENT_USER_GROUP_POLICY_ID (7)
value CERT_SYSTEM_STORE_CURRENT_USER_ID (1)
value CERT_SYSTEM_STORE_DEFER_READ_FLAG (0x20000000)
value CERT_SYSTEM_STORE_LOCAL_MACHINE_ENTERPRISE_ID (9)
value CERT_SYSTEM_STORE_LOCAL_MACHINE_GROUP_POLICY_ID (8)
value CERT_SYSTEM_STORE_LOCAL_MACHINE_ID (2)
value CERT_SYSTEM_STORE_LOCAL_MACHINE_WCOS_ID (10)
value CERT_SYSTEM_STORE_LOCATION_MASK (0x00FF0000)
value CERT_SYSTEM_STORE_LOCATION_SHIFT (16)
value CERT_SYSTEM_STORE_MASK (0xFFFF0000)
value CERT_SYSTEM_STORE_RELOCATE_FLAG (0x80000000)
value CERT_SYSTEM_STORE_SERVICES_ID (5)
value CERT_SYSTEM_STORE_UNPROTECTED_FLAG (0x40000000)
value CERT_SYSTEM_STORE_USERS_ID (6)
value CERT_TIMESTAMP_HASH_USE_TYPE (2)
value CERT_TRUST_AUTO_UPDATE_CA_REVOCATION (0x00000010)
value CERT_TRUST_AUTO_UPDATE_END_REVOCATION (0x00000020)
value CERT_TRUST_BEFORE_DISALLOWED_CA_FILETIME (0x00200000)
value CERT_TRUST_CTL_IS_NOT_SIGNATURE_VALID (0x00040000)
value CERT_TRUST_CTL_IS_NOT_TIME_VALID (0x00020000)
value CERT_TRUST_CTL_IS_NOT_VALID_FOR_USAGE (0x00080000)
value CERT_TRUST_HAS_ALLOW_WEAK_SIGNATURE (0x00020000)
value CERT_TRUST_HAS_AUTO_UPDATE_WEAK_SIGNATURE (0x00008000)
value CERT_TRUST_HAS_CRL_VALIDITY_EXTENDED (0x00001000)
value CERT_TRUST_HAS_EXACT_MATCH_ISSUER (0x00000001)
value CERT_TRUST_HAS_EXCLUDED_NAME_CONSTRAINT (0x00008000)
value CERT_TRUST_HAS_ISSUANCE_CHAIN_POLICY (0x00000200)
value CERT_TRUST_HAS_KEY_MATCH_ISSUER (0x00000002)
value CERT_TRUST_HAS_NAME_MATCH_ISSUER (0x00000004)
value CERT_TRUST_HAS_NOT_DEFINED_NAME_CONSTRAINT (0x00002000)
value CERT_TRUST_HAS_NOT_PERMITTED_NAME_CONSTRAINT (0x00004000)
value CERT_TRUST_HAS_NOT_SUPPORTED_CRITICAL_EXT (0x08000000)
value CERT_TRUST_HAS_NOT_SUPPORTED_NAME_CONSTRAINT (0x00001000)
value CERT_TRUST_HAS_PREFERRED_ISSUER (0x00000100)
value CERT_TRUST_HAS_VALID_NAME_CONSTRAINTS (0x00000400)
value CERT_TRUST_HAS_WEAK_HYGIENE (0x00200000)
value CERT_TRUST_HAS_WEAK_SIGNATURE (0x00100000)
value CERT_TRUST_INVALID_BASIC_CONSTRAINTS (0x00000400)
value CERT_TRUST_INVALID_EXTENSION (0x00000100)
value CERT_TRUST_INVALID_NAME_CONSTRAINTS (0x00000800)
value CERT_TRUST_INVALID_POLICY_CONSTRAINTS (0x00000200)
value CERT_TRUST_IS_CA_TRUSTED (0x00004000)
value CERT_TRUST_IS_COMPLEX_CHAIN (0x00010000)
value CERT_TRUST_IS_CYCLIC (0x00000080)
value CERT_TRUST_IS_EXPLICIT_DISTRUST (0x04000000)
value CERT_TRUST_IS_FROM_EXCLUSIVE_TRUST_STORE (0x00002000)
value CERT_TRUST_IS_KEY_ROLLOVER (0x00000080)
value CERT_TRUST_IS_NOT_SIGNATURE_VALID (0x00000008)
value CERT_TRUST_IS_NOT_TIME_NESTED (0x00000002)
value CERT_TRUST_IS_NOT_TIME_VALID (0x00000001)
value CERT_TRUST_IS_NOT_VALID_FOR_USAGE (0x00000010)
value CERT_TRUST_IS_OFFLINE_REVOCATION (0x01000000)
value CERT_TRUST_IS_PARTIAL_CHAIN (0x00010000)
value CERT_TRUST_IS_PEER_TRUSTED (0x00000800)
value CERT_TRUST_IS_REVOKED (0x00000004)
value CERT_TRUST_IS_SELF_SIGNED (0x00000008)
value CERT_TRUST_IS_UNTRUSTED_ROOT (0x00000020)
value CERT_TRUST_NO_ERROR (0x00000000)
value CERT_TRUST_NO_ISSUANCE_CHAIN_POLICY (0x02000000)
value CERT_TRUST_NO_OCSP_FAILOVER_TO_CRL (0x00000040)
value CERT_TRUST_NO_TIME_CHECK (0x02000000)
value CERT_TRUST_PUB_ALLOW_END_USER_TRUST (0x00000000)
value CERT_TRUST_PUB_ALLOW_ENTERPRISE_ADMIN_TRUST (0x00000002)
value CERT_TRUST_PUB_ALLOW_MACHINE_ADMIN_TRUST (0x00000001)
value CERT_TRUST_PUB_ALLOW_TRUST_MASK (0x00000003)
value CERT_TRUST_PUB_CHECK_PUBLISHER_REV_FLAG (0x00000100)
value CERT_TRUST_PUB_CHECK_TIMESTAMP_REV_FLAG (0x00000200)
value CERT_TRUST_REVOCATION_STATUS_UNKNOWN (0x00000040)
value CERT_TRUST_SSL_HANDSHAKE_OCSP (0x00040000)
value CERT_TRUST_SSL_RECONNECT_OCSP (0x00100000)
value CERT_TRUST_SSL_TIME_VALID (0x01000000)
value CERT_TRUST_SSL_TIME_VALID_OCSP (0x00080000)
value CERT_UNICODE_ATTR_ERR_INDEX_MASK (0x003F)
value CERT_UNICODE_ATTR_ERR_INDEX_SHIFT (16)
value CERT_UNICODE_IS_RDN_ATTRS_FLAG (0x1)
value CERT_UNICODE_RDN_ERR_INDEX_MASK (0x3FF)
value CERT_UNICODE_RDN_ERR_INDEX_SHIFT (22)
value CERT_UNICODE_VALUE_ERR_INDEX_MASK (0x0000FFFF)
value CERT_UNICODE_VALUE_ERR_INDEX_SHIFT (0)
value CERT_VERIFY_ALLOW_MORE_USAGE_FLAG (0x8)
value CERT_VERIFY_CACHE_ONLY_BASED_REVOCATION (0x00000002)
value CERT_VERIFY_INHIBIT_CTL_UPDATE_FLAG (0x1)
value CERT_VERIFY_NO_TIME_CHECK_FLAG (0x4)
value CERT_VERIFY_REV_ACCUMULATIVE_TIMEOUT_FLAG (0x00000004)
value CERT_VERIFY_REV_CHAIN_FLAG (0x00000001)
value CERT_VERIFY_REV_NO_OCSP_FAILOVER_TO_CRL_FLAG (0x00000010)
value CERT_VERIFY_REV_SERVER_OCSP_FLAG (0x00000008)
value CERT_VERIFY_REV_SERVER_OCSP_WIRE_ONLY_FLAG (0x00000020)
value CERT_VERIFY_TRUSTED_SIGNERS_FLAG (0x2)
value CERT_VERIFY_UPDATED_CTL_FLAG (0x1)
value CERT_XML_NAME_STR (4)
value CE_BREAK (0x0010)
value CE_DNS (0x0800)
value CE_FRAME (0x0008)
value CE_IOE (0x0400)
value CE_MODE (0x8000)
value CE_OOP (0x1000)
value CE_OVERRUN (0x0002)
value CE_PTO (0x0200)
value CE_RXOVER (0x0001)
value CE_RXPARITY (0x0004)
value CE_TXFULL (0x0100)
value CFERR_CHOOSEFONTCODES (0x2000)
value CFERR_MAXLESSTHANMIN (0x2002)
value CFERR_NOFONTS (0x2001)
value CFG_CALL_TARGET_CONVERT_EXPORT_SUPPRESSED_TO_VALID ((0x00000004))
value CFG_CALL_TARGET_CONVERT_XFG_TO_CFG ((0x00000010))
value CFG_CALL_TARGET_PROCESSED ((0x00000002))
value CFG_CALL_TARGET_VALID ((0x00000001))
value CFG_CALL_TARGET_VALID_XFG ((0x00000008))
value CFORCEINLINE (FORCEINLINE)
value CFSTR_MIME_NULL (NULL)
value CFS_CANDIDATEPOS (0x0040)
value CFS_DEFAULT (0x0000)
value CFS_EXCLUDE (0x0080)
value CFS_FORCE_POSITION (0x0020)
value CFS_POINT (0x0002)
value CFS_RECT (0x0001)
value CF_ACCEPT (0x0000)
value CF_ANSIONLY (0x00000400L)
value CF_APPLY (0x00000200L)
value CF_BITMAP (2)
value CF_BOTH ((CF_SCREENFONTS | CF_PRINTERFONTS))
value CF_DEFER (0x0002)
value CF_DIB (8)
value CF_DIF (5)
value CF_DSPBITMAP (0x0082)
value CF_DSPENHMETAFILE (0x008E)
value CF_DSPMETAFILEPICT (0x0083)
value CF_DSPTEXT (0x0081)
value CF_EFFECTS (0x00000100L)
value CF_ENABLEHOOK (0x00000008L)
value CF_ENABLETEMPLATE (0x00000010L)
value CF_ENABLETEMPLATEHANDLE (0x00000020L)
value CF_ENHMETAFILE (14)
value CF_FIXEDPITCHONLY (0x00004000L)
value CF_FORCEFONTEXIST (0x00010000L)
value CF_GDIOBJFIRST (0x0300)
value CF_GDIOBJLAST (0x03FF)
value CF_HDROP (15)
value CF_INACTIVEFONTS (0x02000000L)
value CF_INITTOLOGFONTSTRUCT (0x00000040L)
value CF_LIMITSIZE (0x00002000L)
value CF_LOCALE (16)
value CF_MAX (18)
value CF_METAFILEPICT (3)
value CF_NOFACESEL (0x00080000L)
value CF_NOOEMFONTS (CF_NOVECTORFONTS)
value CF_NOSCRIPTSEL (0x00800000L)
value CF_NOSIMULATIONS (0x00001000L)
value CF_NOSIZESEL (0x00200000L)
value CF_NOSTYLESEL (0x00100000L)
value CF_NOVECTORFONTS (0x00000800L)
value CF_NOVERTFONTS (0x01000000L)
value CF_NULL (0)
value CF_OEMTEXT (7)
value CF_OWNERDISPLAY (0x0080)
value CF_PALETTE (9)
value CF_PENDATA (10)
value CF_PRINTERFONTS (0x00000002)
value CF_PRIVATEFIRST (0x0200)
value CF_PRIVATELAST (0x02FF)
value CF_REJECT (0x0001)
value CF_RIFF (11)
value CF_SCALABLEONLY (0x00020000L)
value CF_SCREENFONTS (0x00000001)
value CF_SCRIPTSONLY (CF_ANSIONLY)
value CF_SELECTSCRIPT (0x00400000L)
value CF_SHOWHELP (0x00000004L)
value CF_SYLK (4)
value CF_TEXT (1)
value CF_TIFF (6)
value CF_TTONLY (0x00040000L)
value CF_UNICODETEXT (13)
value CF_USESTYLE (0x00000080L)
value CF_WAVE (12)
value CF_WYSIWYG (0x00008000L)
value CHANGER_BAR_CODE_SCANNER_INSTALLED (0x00000001)
value CHANGER_CARTRIDGE_MAGAZINE (0x00000100)
value CHANGER_CLEANER_ACCESS_NOT_VALID (0x00040000)
value CHANGER_CLEANER_AUTODISMOUNT (0x80000004)
value CHANGER_CLEANER_OPS_NOT_SUPPORTED (0x80000040)
value CHANGER_CLEANER_SLOT (0x00000040)
value CHANGER_CLOSE_IEPORT (0x00000004)
value CHANGER_DEVICE_REINITIALIZE_CAPABLE (0x08000000)
value CHANGER_DRIVE_CLEANING_REQUIRED (0x00010000)
value CHANGER_DRIVE_EMPTY_ON_DOOR_ACCESS (0x20000000)
value CHANGER_EXCHANGE_MEDIA (0x00000020)
value CHANGER_IEPORT_USER_CONTROL_CLOSE (0x80000100)
value CHANGER_IEPORT_USER_CONTROL_OPEN (0x80000080)
value CHANGER_INIT_ELEM_STAT_WITH_RANGE (0x00000002)
value CHANGER_KEYPAD_ENABLE_DISABLE (0x10000000)
value CHANGER_LOCK_UNLOCK (0x00000080)
value CHANGER_MEDIUM_FLIP (0x00000200)
value CHANGER_MOVE_EXTENDS_IEPORT (0x80000200)
value CHANGER_MOVE_RETRACTS_IEPORT (0x80000400)
value CHANGER_OPEN_IEPORT (0x00000008)
value CHANGER_POSITION_TO_ELEMENT (0x00000400)
value CHANGER_PREDISMOUNT_ALIGN_TO_DRIVE (0x80000002)
value CHANGER_PREDISMOUNT_ALIGN_TO_SLOT (0x80000001)
value CHANGER_PREDISMOUNT_EJECT_REQUIRED (0x00020000)
value CHANGER_PREMOUNT_EJECT_REQUIRED (0x00080000)
value CHANGER_REPORT_IEPORT_STATE (0x00000800)
value CHANGER_RESERVED_BIT (0x80000000)
value CHANGER_RTN_MEDIA_TO_ORIGINAL_ADDR (0x80000020)
value CHANGER_SERIAL_NUMBER_VALID (0x04000000)
value CHANGER_SLOTS_USE_TRAYS (0x80000010)
value CHANGER_STATUS_NON_VOLATILE (0x00000010)
value CHANGER_STORAGE_DRIVE (0x00001000)
value CHANGER_STORAGE_IEPORT (0x00002000)
value CHANGER_STORAGE_SLOT (0x00004000)
value CHANGER_STORAGE_TRANSPORT (0x00008000)
value CHANGER_TO_DRIVE (0x08)
value CHANGER_TO_IEPORT (0x04)
value CHANGER_TO_SLOT (0x02)
value CHANGER_TO_TRANSPORT (0x01)
value CHANGER_TRUE_EXCHANGE_CAPABLE (0x80000008)
value CHANGER_VOLUME_ASSERT (0x00400000)
value CHANGER_VOLUME_IDENTIFICATION (0x00100000)
value CHANGER_VOLUME_REPLACE (0x00800000)
value CHANGER_VOLUME_SEARCH (0x00200000)
value CHANGER_VOLUME_UNDEFINE (0x01000000)
value CHAR_BIT (8)
value CHAR_MAX (SCHAR_MAX)
value CHAR_MIN (SCHAR_MIN)
value CHECKJPEGFORMAT (4119)
value CHECKPNGFORMAT (4120)
value CHECKSUM_TYPE_ECC ((3))
value CHECKSUM_TYPE_FIRST_UNUSED_TYPE ((4))
value CHECKSUM_TYPE_NONE ((0))
value CHECKSUM_TYPE_UNCHANGED ((-1))
value CHILDID_SELF (0)
value CLAIM_SECURITY_ATTRIBUTES_INFORMATION_VERSION (CLAIM_SECURITY_ATTRIBUTES_INFORMATION_VERSION_V1)
value CLAIM_SECURITY_ATTRIBUTE_CUSTOM_FLAGS (0xFFFF0000)
value CLAIM_SECURITY_ATTRIBUTE_DISABLED (0x0010)
value CLAIM_SECURITY_ATTRIBUTE_DISABLED_BY_DEFAULT (0x0008)
value CLAIM_SECURITY_ATTRIBUTE_MANDATORY (0x0020)
value CLAIM_SECURITY_ATTRIBUTE_NON_INHERITABLE (0x0001)
value CLAIM_SECURITY_ATTRIBUTE_TYPE_BOOLEAN (0x06)
value CLAIM_SECURITY_ATTRIBUTE_TYPE_FQBN (0x04)
value CLAIM_SECURITY_ATTRIBUTE_TYPE_INVALID (0x00)
value CLAIM_SECURITY_ATTRIBUTE_TYPE_OCTET_STRING (0x10)
value CLAIM_SECURITY_ATTRIBUTE_TYPE_SID (0x05)
value CLAIM_SECURITY_ATTRIBUTE_TYPE_STRING (0x03)
value CLAIM_SECURITY_ATTRIBUTE_USE_FOR_DENY_ONLY (0x0004)
value CLAIM_SECURITY_ATTRIBUTE_VALID_FLAGS (( CLAIM_SECURITY_ATTRIBUTE_NON_INHERITABLE | CLAIM_SECURITY_ATTRIBUTE_VALUE_CASE_SENSITIVE | CLAIM_SECURITY_ATTRIBUTE_USE_FOR_DENY_ONLY | CLAIM_SECURITY_ATTRIBUTE_DISABLED_BY_DEFAULT | CLAIM_SECURITY_ATTRIBUTE_DISABLED | CLAIM_SECURITY_ATTRIBUTE_MANDATORY ))
value CLAIM_SECURITY_ATTRIBUTE_VALUE_CASE_SENSITIVE (0x0002)
value CLASSFACTORY_E_FIRST (0x80040110L)
value CLASSFACTORY_E_LAST (0x8004011FL)
value CLASSFACTORY_S_FIRST (0x00040110L)
value CLASSFACTORY_S_LAST (0x0004011FL)
value CLASS_E_CLASSNOTAVAILABLE (_HRESULT_TYPEDEF_(0x80040111L))
value CLASS_E_NOAGGREGATION (_HRESULT_TYPEDEF_(0x80040110L))
value CLASS_E_NOTLICENSED (_HRESULT_TYPEDEF_(0x80040112L))
value CLEARTYPE_NATURAL_QUALITY (6)
value CLEARTYPE_QUALITY (5)
value CLIENTSITE_E_FIRST (0x80040190L)
value CLIENTSITE_E_LAST (0x8004019FL)
value CLIENTSITE_S_FIRST (0x00040190L)
value CLIENTSITE_S_LAST (0x0004019FL)
value CLIPBRD_E_BAD_DATA (_HRESULT_TYPEDEF_(0x800401D3L))
value CLIPBRD_E_CANT_CLOSE (_HRESULT_TYPEDEF_(0x800401D4L))
value CLIPBRD_E_CANT_EMPTY (_HRESULT_TYPEDEF_(0x800401D1L))
value CLIPBRD_E_CANT_OPEN (_HRESULT_TYPEDEF_(0x800401D0L))
value CLIPBRD_E_CANT_SET (_HRESULT_TYPEDEF_(0x800401D2L))
value CLIPBRD_E_FIRST (0x800401D0L)
value CLIPBRD_E_LAST (0x800401DFL)
value CLIPBRD_S_FIRST (0x000401D0L)
value CLIPBRD_S_LAST (0x000401DFL)
value CLIPCAPS (36)
value CLIP_CHARACTER_PRECIS (1)
value CLIP_DEFAULT_PRECIS (0)
value CLIP_MASK (0xf)
value CLIP_STROKE_PRECIS (2)
value CLIP_TO_PATH (4097)
value CLK_TCK (CLOCKS_PER_SEC)
value CLOSECHANNEL (4112)
value CLRBREAK (9)
value CLRDTR (6)
value CLRRTS (4)
value CLR_INVALID (0xFFFFFFFF)
value CLSCTX_ALL ((CLSCTX_INPROC_SERVER| CLSCTX_INPROC_HANDLER| CLSCTX_LOCAL_SERVER| CLSCTX_REMOTE_SERVER))
value CLSCTX_INPROC ((CLSCTX_INPROC_SERVER|CLSCTX_INPROC_HANDLER))
value CLSCTX_SERVER ((CLSCTX_INPROC_SERVER|CLSCTX_LOCAL_SERVER|CLSCTX_REMOTE_SERVER))
value CLSCTX_VALID_MASK ((CLSCTX_INPROC_SERVER | CLSCTX_INPROC_HANDLER | CLSCTX_LOCAL_SERVER | CLSCTX_INPROC_SERVER16 | CLSCTX_REMOTE_SERVER | CLSCTX_NO_CODE_DOWNLOAD | CLSCTX_NO_CUSTOM_MARSHAL | CLSCTX_ENABLE_CODE_DOWNLOAD | CLSCTX_NO_FAILURE_LOG | CLSCTX_DISABLE_AAA | CLSCTX_ENABLE_AAA | CLSCTX_FROM_DEFAULT_CONTEXT | CLSCTX_ACTIVATE_X86_SERVER | CLSCTX_ACTIVATE_64_BIT_SERVER | CLSCTX_ENABLE_CLOAKING | CLSCTX_APPCONTAINER | CLSCTX_ACTIVATE_AAA_AS_IU | CLSCTX_RESERVED6 | CLSCTX_ACTIVATE_ARM32_SERVER | CLSCTX_ALLOW_LOWER_TRUST_REGISTRATION | CLSCTX_PS_DLL))
value CLSID_NULL (GUID_NULL)
value CMAPI (DECLSPEC_IMPORT)
value CMC_ADD_ATTRIBUTES (((LPCSTR) 63))
value CMC_ADD_EXTENSIONS (((LPCSTR) 62))
value CMC_DATA (((LPCSTR) 59))
value CMC_FAIL_BAD_ALG (0)
value CMC_FAIL_BAD_CERT_ID (4)
value CMC_FAIL_BAD_IDENTITY (7)
value CMC_FAIL_BAD_MESSAGE_CHECK (1)
value CMC_FAIL_BAD_REQUEST (2)
value CMC_FAIL_BAD_TIME (3)
value CMC_FAIL_INTERNAL_CA_ERROR (11)
value CMC_FAIL_MUST_ARCHIVE_KEYS (6)
value CMC_FAIL_NO_KEY_REUSE (10)
value CMC_FAIL_POP_FAILED (9)
value CMC_FAIL_POP_REQUIRED (8)
value CMC_FAIL_TRY_LATER (12)
value CMC_FAIL_UNSUPORTED_EXT (5)
value CMC_OTHER_INFO_FAIL_CHOICE (1)
value CMC_OTHER_INFO_NO_CHOICE (0)
value CMC_OTHER_INFO_PEND_CHOICE (2)
value CMC_RESPONSE (((LPCSTR) 60))
value CMC_STATUS (((LPCSTR) 61))
value CMC_STATUS_CONFIRM_REQUIRED (5)
value CMC_STATUS_FAILED (2)
value CMC_STATUS_NO_SUPPORT (4)
value CMC_STATUS_PENDING (3)
value CMC_STATUS_SUCCESS (0)
value CMC_TAGGED_CERT_REQUEST_CHOICE (1)
value CMSGDATA_ALIGN (WSA_CMSGDATA_ALIGN)
value CMSGHDR_ALIGN (WSA_CMSGHDR_ALIGN)
value CMSG_ATTR_CERT_COUNT_PARAM (31)
value CMSG_ATTR_CERT_PARAM (32)
value CMSG_AUTHENTICATED_ATTRIBUTES_FLAG (0x00000008)
value CMSG_BARE_CONTENT_FLAG (0x00000001)
value CMSG_BARE_CONTENT_PARAM (3)
value CMSG_CERT_COUNT_PARAM (11)
value CMSG_CERT_PARAM (12)
value CMSG_CMS_ENCAPSULATED_CONTENT_FLAG (0x00000040)
value CMSG_CMS_ENCAPSULATED_CTL_FLAG (0x00008000)
value CMSG_CMS_RECIPIENT_COUNT_PARAM (33)
value CMSG_CMS_RECIPIENT_ENCRYPTED_KEY_INDEX_PARAM (35)
value CMSG_CMS_RECIPIENT_INDEX_PARAM (34)
value CMSG_CMS_RECIPIENT_INFO_PARAM (36)
value CMSG_CMS_SIGNER_INFO_PARAM (39)
value CMSG_COMPUTED_HASH_PARAM (22)
value CMSG_CONTENTS_OCTETS_FLAG (0x00000010)
value CMSG_CONTENT_ENCRYPT_FREE_OBJID_FLAG (0x00000002)
value CMSG_CONTENT_ENCRYPT_FREE_PARA_FLAG (0x00000001)
value CMSG_CONTENT_ENCRYPT_PAD_ENCODED_LEN_FLAG (0x00000001)
value CMSG_CONTENT_ENCRYPT_RELEASE_CONTEXT_FLAG (0x00008000)
value CMSG_CONTENT_PARAM (2)
value CMSG_CRL_COUNT_PARAM (13)
value CMSG_CRL_PARAM (14)
value CMSG_CRYPT_RELEASE_CONTEXT_FLAG (0x00008000)
value CMSG_CTRL_ADD_ATTR_CERT (14)
value CMSG_CTRL_ADD_CERT (10)
value CMSG_CTRL_ADD_CMS_SIGNER_INFO (20)
value CMSG_CTRL_ADD_CRL (12)
value CMSG_CTRL_ADD_SIGNER (6)
value CMSG_CTRL_ADD_SIGNER_UNAUTH_ATTR (8)
value CMSG_CTRL_DECRYPT (2)
value CMSG_CTRL_DEL_ATTR_CERT (15)
value CMSG_CTRL_DEL_CERT (11)
value CMSG_CTRL_DEL_CRL (13)
value CMSG_CTRL_DEL_SIGNER (7)
value CMSG_CTRL_DEL_SIGNER_UNAUTH_ATTR (9)
value CMSG_CTRL_ENABLE_STRONG_SIGNATURE (21)
value CMSG_CTRL_KEY_AGREE_DECRYPT (17)
value CMSG_CTRL_KEY_TRANS_DECRYPT (16)
value CMSG_CTRL_MAIL_LIST_DECRYPT (18)
value CMSG_CTRL_VERIFY_HASH (5)
value CMSG_CTRL_VERIFY_SIGNATURE (1)
value CMSG_CTRL_VERIFY_SIGNATURE_EX (19)
value CMSG_DATA (1)
value CMSG_DEFAULT_INSTALLABLE_FUNC_OID (((LPCSTR) 1))
value CMSG_DETACHED_FLAG (0x00000004)
value CMSG_ENCODED_MESSAGE (29)
value CMSG_ENCODED_SIGNER (28)
value CMSG_ENCODE_HASHED_SUBJECT_IDENTIFIER_FLAG (0x2)
value CMSG_ENCODE_SORTED_CTL_FLAG (0x1)
value CMSG_ENCODING_TYPE_MASK (0xFFFF0000)
value CMSG_ENCRYPTED (6)
value CMSG_ENCRYPTED_DIGEST (27)
value CMSG_ENCRYPT_PARAM (26)
value CMSG_ENVELOPED (3)
value CMSG_ENVELOPED_DATA_CMS_VERSION (CMSG_ENVELOPED_DATA_V2)
value CMSG_ENVELOPE_ALGORITHM_PARAM (15)
value CMSG_FIRSTHDR (WSA_CMSG_FIRSTHDR)
value CMSG_HASHED (5)
value CMSG_HASHED_DATA_CMS_VERSION (CMSG_HASHED_DATA_V2)
value CMSG_HASH_ALGORITHM_PARAM (20)
value CMSG_HASH_DATA_PARAM (21)
value CMSG_INDEFINITE_LENGTH ((0xFFFFFFFF))
value CMSG_INNER_CONTENT_TYPE_PARAM (4)
value CMSG_KEY_AGREE_ENCRYPT_FREE_MATERIAL_FLAG (0x00000002)
value CMSG_KEY_AGREE_ENCRYPT_FREE_OBJID_FLAG (0x00000020)
value CMSG_KEY_AGREE_ENCRYPT_FREE_PARA_FLAG (0x00000001)
value CMSG_KEY_AGREE_ENCRYPT_FREE_PUBKEY_ALG_FLAG (0x00000004)
value CMSG_KEY_AGREE_ENCRYPT_FREE_PUBKEY_BITS_FLAG (0x00000010)
value CMSG_KEY_AGREE_ENCRYPT_FREE_PUBKEY_PARA_FLAG (0x00000008)
value CMSG_KEY_AGREE_EPHEMERAL_KEY_CHOICE (1)
value CMSG_KEY_AGREE_ORIGINATOR_CERT (1)
value CMSG_KEY_AGREE_ORIGINATOR_PUBLIC_KEY (2)
value CMSG_KEY_AGREE_RECIPIENT (2)
value CMSG_KEY_AGREE_STATIC_KEY_CHOICE (2)
value CMSG_KEY_AGREE_VERSION (CMSG_ENVELOPED_RECIPIENT_V3)
value CMSG_KEY_TRANS_CMS_VERSION (CMSG_ENVELOPED_RECIPIENT_V2)
value CMSG_KEY_TRANS_ENCRYPT_FREE_OBJID_FLAG (0x00000002)
value CMSG_KEY_TRANS_ENCRYPT_FREE_PARA_FLAG (0x00000001)
value CMSG_KEY_TRANS_RECIPIENT (1)
value CMSG_LEN (WSA_CMSG_LEN)
value CMSG_LENGTH_ONLY_FLAG (0x00000002)
value CMSG_MAIL_LIST_ENCRYPT_FREE_OBJID_FLAG (0x00000002)
value CMSG_MAIL_LIST_ENCRYPT_FREE_PARA_FLAG (0x00000001)
value CMSG_MAIL_LIST_HANDLE_KEY_CHOICE (1)
value CMSG_MAIL_LIST_RECIPIENT (3)
value CMSG_MAIL_LIST_VERSION (CMSG_ENVELOPED_RECIPIENT_V4)
value CMSG_MAX_LENGTH_FLAG (0x00000020)
value CMSG_NXTHDR (WSA_CMSG_NXTHDR)
value CMSG_RECIPIENT_COUNT_PARAM (17)
value CMSG_RECIPIENT_INDEX_PARAM (18)
value CMSG_RECIPIENT_INFO_PARAM (19)
value CMSG_SIGNED (2)
value CMSG_SIGNED_AND_ENVELOPED (4)
value CMSG_SIGNED_DATA_CMS_VERSION (CMSG_SIGNED_DATA_V3)
value CMSG_SIGNED_DATA_NO_SIGN_FLAG (0x00000080)
value CMSG_SIGNER_AUTH_ATTR_PARAM (9)
value CMSG_SIGNER_CERT_ID_PARAM (38)
value CMSG_SIGNER_CERT_INFO_PARAM (7)
value CMSG_SIGNER_COUNT_PARAM (5)
value CMSG_SIGNER_HASH_ALGORITHM_PARAM (8)
value CMSG_SIGNER_INFO_CMS_VERSION (CMSG_SIGNER_INFO_V3)
value CMSG_SIGNER_INFO_PARAM (6)
value CMSG_SIGNER_ONLY_FLAG (0x2)
value CMSG_SIGNER_UNAUTH_ATTR_PARAM (10)
value CMSG_SPACE (WSA_CMSG_SPACE)
value CMSG_TRUSTED_SIGNER_FLAG (0x1)
value CMSG_TYPE_PARAM (1)
value CMSG_UNPROTECTED_ATTR_PARAM (37)
value CMSG_USE_SIGNER_INDEX_FLAG (0x4)
value CMSG_VERIFY_COUNTER_SIGN_ENABLE_STRONG_FLAG (0x00000001)
value CMSG_VERIFY_SIGNER_CERT (2)
value CMSG_VERIFY_SIGNER_CHAIN (3)
value CMSG_VERIFY_SIGNER_NULL (4)
value CMSG_VERIFY_SIGNER_PUBKEY (1)
value CMSG_VERSION_PARAM (30)
value CMS_SIGNER_INFO (((LPCSTR) 501))
value CM_CMYK_COLOR (0x00000004)
value CM_DEVICE_ICM (0x00000001)
value CM_GAMMA_RAMP (0x00000002)
value CM_IN_GAMUT (0)
value CM_NONE (0x00000000)
value CM_OUT_OF_GAMUT (255)
value CM_SERVICE_MEASURED_BOOT_LOAD (0x00000020)
value CM_SERVICE_NETWORK_BOOT_LOAD (0x00000001)
value CM_SERVICE_RAM_DISK_BOOT_LOAD (0x00000100)
value CM_SERVICE_SD_DISK_BOOT_LOAD (0x00000008)
value CM_SERVICE_USB_DISK_BOOT_LOAD (0x00000004)
value CM_SERVICE_VALID_PROMOTION_MASK ((CM_SERVICE_NETWORK_BOOT_LOAD | CM_SERVICE_VIRTUAL_DISK_BOOT_LOAD | CM_SERVICE_USB_DISK_BOOT_LOAD | CM_SERVICE_SD_DISK_BOOT_LOAD | CM_SERVICE_USB3_DISK_BOOT_LOAD | CM_SERVICE_MEASURED_BOOT_LOAD | CM_SERVICE_VERIFIER_BOOT_LOAD | CM_SERVICE_WINPE_BOOT_LOAD | CM_SERVICE_RAM_DISK_BOOT_LOAD))
value CM_SERVICE_VERIFIER_BOOT_LOAD (0x00000040)
value CM_SERVICE_VIRTUAL_DISK_BOOT_LOAD (0x00000002)
value CM_SERVICE_WINPE_BOOT_LOAD (0x00000080)
value CNG_RSA_PRIVATE_KEY_BLOB (((LPCSTR) 83))
value CNG_RSA_PUBLIC_KEY_BLOB (((LPCSTR) 72))
value CODEPAGE_ENUMPROC (CODEPAGE_ENUMPROCA)
value COLORMATCHTOTARGET_EMBEDED (0x00000001)
value COLORMGMTCAPS (121)
value COLORMGMTDLGORD (1551)
value COLOROKSTRING (COLOROKSTRINGA)
value COLORONCOLOR (3)
value COLORRES (108)
value COLOR_ACTIVEBORDER (10)
value COLOR_ACTIVECAPTION (2)
value COLOR_ADJ_MAX ((SHORT)100)
value COLOR_ADJ_MIN ((SHORT)-100)
value COLOR_APPWORKSPACE (12)
value COLOR_BACKGROUND (1)
value COLOR_BTNFACE (15)
value COLOR_BTNHIGHLIGHT (20)
value COLOR_BTNHILIGHT (COLOR_BTNHIGHLIGHT)
value COLOR_BTNSHADOW (16)
value COLOR_BTNTEXT (18)
value COLOR_CAPTIONTEXT (9)
value COLOR_DESKTOP (COLOR_BACKGROUND)
value COLOR_GRADIENTACTIVECAPTION (27)
value COLOR_GRADIENTINACTIVECAPTION (28)
value COLOR_GRAYTEXT (17)
value COLOR_HIGHLIGHT (13)
value COLOR_HIGHLIGHTTEXT (14)
value COLOR_HOTLIGHT (26)
value COLOR_INACTIVEBORDER (11)
value COLOR_INACTIVECAPTION (3)
value COLOR_INACTIVECAPTIONTEXT (19)
value COLOR_INFOBK (24)
value COLOR_INFOTEXT (23)
value COLOR_MENU (4)
value COLOR_MENUBAR (30)
value COLOR_MENUHILIGHT (29)
value COLOR_MENUTEXT (7)
value COLOR_SCROLLBAR (0)
value COLOR_WINDOW (5)
value COLOR_WINDOWFRAME (6)
value COLOR_WINDOWTEXT (8)
value COMADMIN_E_ALREADYINSTALLED (_HRESULT_TYPEDEF_(0x80110404L))
value COMADMIN_E_AMBIGUOUS_APPLICATION_NAME (_HRESULT_TYPEDEF_(0x8011045CL))
value COMADMIN_E_AMBIGUOUS_PARTITION_NAME (_HRESULT_TYPEDEF_(0x8011045DL))
value COMADMIN_E_APPDIRNOTFOUND (_HRESULT_TYPEDEF_(0x8011041FL))
value COMADMIN_E_APPLICATIONEXISTS (_HRESULT_TYPEDEF_(0x8011040BL))
value COMADMIN_E_APPLID_MATCHES_CLSID (_HRESULT_TYPEDEF_(0x80110446L))
value COMADMIN_E_APP_FILE_READFAIL (_HRESULT_TYPEDEF_(0x80110408L))
value COMADMIN_E_APP_FILE_VERSION (_HRESULT_TYPEDEF_(0x80110409L))
value COMADMIN_E_APP_FILE_WRITEFAIL (_HRESULT_TYPEDEF_(0x80110407L))
value COMADMIN_E_APP_NOT_RUNNING (_HRESULT_TYPEDEF_(0x8011080AL))
value COMADMIN_E_AUTHENTICATIONLEVEL (_HRESULT_TYPEDEF_(0x80110413L))
value COMADMIN_E_BADPATH (_HRESULT_TYPEDEF_(0x8011040AL))
value COMADMIN_E_BADREGISTRYLIBID (_HRESULT_TYPEDEF_(0x8011041EL))
value COMADMIN_E_BADREGISTRYPROGID (_HRESULT_TYPEDEF_(0x80110412L))
value COMADMIN_E_BASEPARTITION_REQUIRED_IN_SET (_HRESULT_TYPEDEF_(0x8011081FL))
value COMADMIN_E_BASE_PARTITION_ONLY (_HRESULT_TYPEDEF_(0x80110450L))
value COMADMIN_E_CANNOT_ALIAS_EVENTCLASS (_HRESULT_TYPEDEF_(0x80110820L))
value COMADMIN_E_CANTCOPYFILE (_HRESULT_TYPEDEF_(0x8011040DL))
value COMADMIN_E_CANTMAKEINPROCSERVICE (_HRESULT_TYPEDEF_(0x80110814L))
value COMADMIN_E_CANTRECYCLELIBRARYAPPS (_HRESULT_TYPEDEF_(0x8011080FL))
value COMADMIN_E_CANTRECYCLESERVICEAPPS (_HRESULT_TYPEDEF_(0x80110811L))
value COMADMIN_E_CANT_SUBSCRIBE_TO_COMPONENT (_HRESULT_TYPEDEF_(0x8011044DL))
value COMADMIN_E_CAN_NOT_EXPORT_APP_PROXY (_HRESULT_TYPEDEF_(0x8011044AL))
value COMADMIN_E_CAN_NOT_EXPORT_SYS_APP (_HRESULT_TYPEDEF_(0x8011044CL))
value COMADMIN_E_CAN_NOT_START_APP (_HRESULT_TYPEDEF_(0x8011044BL))
value COMADMIN_E_CAT_BITNESSMISMATCH (_HRESULT_TYPEDEF_(0x80110482L))
value COMADMIN_E_CAT_DUPLICATE_PARTITION_NAME (_HRESULT_TYPEDEF_(0x80110457L))
value COMADMIN_E_CAT_IMPORTED_COMPONENTS_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x8011045BL))
value COMADMIN_E_CAT_INVALID_PARTITION_NAME (_HRESULT_TYPEDEF_(0x80110458L))
value COMADMIN_E_CAT_PARTITION_IN_USE (_HRESULT_TYPEDEF_(0x80110459L))
value COMADMIN_E_CAT_PAUSE_RESUME_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80110485L))
value COMADMIN_E_CAT_SERVERFAULT (_HRESULT_TYPEDEF_(0x80110486L))
value COMADMIN_E_CAT_UNACCEPTABLEBITNESS (_HRESULT_TYPEDEF_(0x80110483L))
value COMADMIN_E_CAT_WRONGAPPBITNESS (_HRESULT_TYPEDEF_(0x80110484L))
value COMADMIN_E_CLSIDORIIDMISMATCH (_HRESULT_TYPEDEF_(0x80110418L))
value COMADMIN_E_COMPFILE_BADTLB (_HRESULT_TYPEDEF_(0x80110428L))
value COMADMIN_E_COMPFILE_CLASSNOTAVAIL (_HRESULT_TYPEDEF_(0x80110427L))
value COMADMIN_E_COMPFILE_DOESNOTEXIST (_HRESULT_TYPEDEF_(0x80110424L))
value COMADMIN_E_COMPFILE_GETCLASSOBJ (_HRESULT_TYPEDEF_(0x80110426L))
value COMADMIN_E_COMPFILE_LOADDLLFAIL (_HRESULT_TYPEDEF_(0x80110425L))
value COMADMIN_E_COMPFILE_NOREGISTRAR (_HRESULT_TYPEDEF_(0x80110434L))
value COMADMIN_E_COMPFILE_NOTINSTALLABLE (_HRESULT_TYPEDEF_(0x80110429L))
value COMADMIN_E_COMPONENTEXISTS (_HRESULT_TYPEDEF_(0x80110439L))
value COMADMIN_E_COMP_MOVE_BAD_DEST (_HRESULT_TYPEDEF_(0x8011042EL))
value COMADMIN_E_COMP_MOVE_DEST (_HRESULT_TYPEDEF_(0x8011081DL))
value COMADMIN_E_COMP_MOVE_LOCKED (_HRESULT_TYPEDEF_(0x8011042DL))
value COMADMIN_E_COMP_MOVE_PRIVATE (_HRESULT_TYPEDEF_(0x8011081EL))
value COMADMIN_E_COMP_MOVE_SOURCE (_HRESULT_TYPEDEF_(0x8011081CL))
value COMADMIN_E_COREQCOMPINSTALLED (_HRESULT_TYPEDEF_(0x80110435L))
value COMADMIN_E_DEFAULT_PARTITION_NOT_IN_SET (_HRESULT_TYPEDEF_(0x80110816L))
value COMADMIN_E_DLLLOADFAILED (_HRESULT_TYPEDEF_(0x8011041DL))
value COMADMIN_E_DLLREGISTERSERVER (_HRESULT_TYPEDEF_(0x8011041AL))
value COMADMIN_E_EVENTCLASS_CANT_BE_SUBSCRIBER (_HRESULT_TYPEDEF_(0x8011044EL))
value COMADMIN_E_FILE_PARTITION_DUPLICATE_FILES (_HRESULT_TYPEDEF_(0x8011045AL))
value COMADMIN_E_INVALIDUSERIDS (_HRESULT_TYPEDEF_(0x80110410L))
value COMADMIN_E_INVALID_PARTITION (_HRESULT_TYPEDEF_(0x8011080BL))
value COMADMIN_E_KEYMISSING (_HRESULT_TYPEDEF_(0x80110403L))
value COMADMIN_E_LEGACYCOMPS_NOT_ALLOWED_IN_NONBASE_PARTITIONS (_HRESULT_TYPEDEF_(0x8011081BL))
value COMADMIN_E_LIB_APP_PROXY_INCOMPATIBLE (_HRESULT_TYPEDEF_(0x8011044FL))
value COMADMIN_E_MIG_SCHEMANOTFOUND (_HRESULT_TYPEDEF_(0x80110481L))
value COMADMIN_E_MIG_VERSIONNOTSUPPORTED (_HRESULT_TYPEDEF_(0x80110480L))
value COMADMIN_E_NOREGISTRYCLSID (_HRESULT_TYPEDEF_(0x80110411L))
value COMADMIN_E_NOSERVERSHARE (_HRESULT_TYPEDEF_(0x8011041BL))
value COMADMIN_E_NOTCHANGEABLE (_HRESULT_TYPEDEF_(0x8011042AL))
value COMADMIN_E_NOTDELETEABLE (_HRESULT_TYPEDEF_(0x8011042BL))
value COMADMIN_E_NOTINREGISTRY (_HRESULT_TYPEDEF_(0x8011043EL))
value COMADMIN_E_NOUSER (_HRESULT_TYPEDEF_(0x8011040FL))
value COMADMIN_E_OBJECTERRORS (_HRESULT_TYPEDEF_(0x80110401L))
value COMADMIN_E_OBJECTEXISTS (_HRESULT_TYPEDEF_(0x80110438L))
value COMADMIN_E_OBJECTINVALID (_HRESULT_TYPEDEF_(0x80110402L))
value COMADMIN_E_OBJECTNOTPOOLABLE (_HRESULT_TYPEDEF_(0x8011043FL))
value COMADMIN_E_OBJECT_DOES_NOT_EXIST (_HRESULT_TYPEDEF_(0x80110809L))
value COMADMIN_E_OBJECT_PARENT_MISSING (_HRESULT_TYPEDEF_(0x80110808L))
value COMADMIN_E_PARTITIONS_DISABLED (_HRESULT_TYPEDEF_(0x80110824L))
value COMADMIN_E_PARTITION_ACCESSDENIED (_HRESULT_TYPEDEF_(0x80110818L))
value COMADMIN_E_PARTITION_MSI_ONLY (_HRESULT_TYPEDEF_(0x80110819L))
value COMADMIN_E_PAUSEDPROCESSMAYNOTBERECYCLED (_HRESULT_TYPEDEF_(0x80110813L))
value COMADMIN_E_PRIVATE_ACCESSDENIED (_HRESULT_TYPEDEF_(0x80110821L))
value COMADMIN_E_PROCESSALREADYRECYCLED (_HRESULT_TYPEDEF_(0x80110812L))
value COMADMIN_E_PROGIDINUSEBYCLSID (_HRESULT_TYPEDEF_(0x80110815L))
value COMADMIN_E_PROPERTYSAVEFAILED (_HRESULT_TYPEDEF_(0x80110437L))
value COMADMIN_E_PROPERTY_OVERFLOW (_HRESULT_TYPEDEF_(0x8011043CL))
value COMADMIN_E_RECYCLEDPROCESSMAYNOTBEPAUSED (_HRESULT_TYPEDEF_(0x80110817L))
value COMADMIN_E_REGDB_ALREADYRUNNING (_HRESULT_TYPEDEF_(0x80110475L))
value COMADMIN_E_REGDB_NOTINITIALIZED (_HRESULT_TYPEDEF_(0x80110472L))
value COMADMIN_E_REGDB_NOTOPEN (_HRESULT_TYPEDEF_(0x80110473L))
value COMADMIN_E_REGDB_SYSTEMERR (_HRESULT_TYPEDEF_(0x80110474L))
value COMADMIN_E_REGFILE_CORRUPT (_HRESULT_TYPEDEF_(0x8011043BL))
value COMADMIN_E_REGISTERTLB (_HRESULT_TYPEDEF_(0x80110430L))
value COMADMIN_E_REGISTRARFAILED (_HRESULT_TYPEDEF_(0x80110423L))
value COMADMIN_E_REGISTRY_ACCESSDENIED (_HRESULT_TYPEDEF_(0x80110823L))
value COMADMIN_E_REMOTEINTERFACE (_HRESULT_TYPEDEF_(0x80110419L))
value COMADMIN_E_REQUIRES_DIFFERENT_PLATFORM (_HRESULT_TYPEDEF_(0x80110449L))
value COMADMIN_E_ROLEEXISTS (_HRESULT_TYPEDEF_(0x8011040CL))
value COMADMIN_E_ROLE_DOES_NOT_EXIST (_HRESULT_TYPEDEF_(0x80110447L))
value COMADMIN_E_SAFERINVALID (_HRESULT_TYPEDEF_(0x80110822L))
value COMADMIN_E_SERVICENOTINSTALLED (_HRESULT_TYPEDEF_(0x80110436L))
value COMADMIN_E_SESSION (_HRESULT_TYPEDEF_(0x8011042CL))
value COMADMIN_E_START_APP_DISABLED (_HRESULT_TYPEDEF_(0x80110451L))
value COMADMIN_E_START_APP_NEEDS_COMPONENTS (_HRESULT_TYPEDEF_(0x80110448L))
value COMADMIN_E_SVCAPP_NOT_POOLABLE_OR_RECYCLABLE (_HRESULT_TYPEDEF_(0x8011080DL))
value COMADMIN_E_SYSTEMAPP (_HRESULT_TYPEDEF_(0x80110433L))
value COMADMIN_E_USERPASSWDNOTVALID (_HRESULT_TYPEDEF_(0x80110414L))
value COMADMIN_E_USER_IN_SET (_HRESULT_TYPEDEF_(0x8011080EL))
value COMMON_LVB_GRID_HORIZONTAL (0x0400)
value COMMON_LVB_GRID_LVERTICAL (0x0800)
value COMMON_LVB_GRID_RVERTICAL (0x1000)
value COMMON_LVB_LEADING_BYTE (0x0100)
value COMMON_LVB_REVERSE_VIDEO (0x4000)
value COMMON_LVB_SBCSDBCS (0x0300)
value COMMON_LVB_TRAILING_BYTE (0x0200)
value COMMON_LVB_UNDERSCORE (0x8000)
value COMMPROP_INITIALIZED (((DWORD)0xE73CF52E))
value COMPLEXREGION (3)
value COMPONENT_KTM (0x01)
value COMPONENT_VALID_FLAGS ((COMPONENT_KTM))
value COMPRESSION_ENGINE_HIBER ((0x0200))
value COMPRESSION_ENGINE_MAXIMUM ((0x0100))
value COMPRESSION_ENGINE_STANDARD ((0x0000))
value COMPRESSION_FORMAT_DEFAULT ((0x0001))
value COMPRESSION_FORMAT_NONE ((0x0000))
value COMPRESSION_FORMAT_XPRESS ((0x0003))
value COMPRESSION_FORMAT_XPRESS_HUFF ((0x0004))
value COMQC_E_APPLICATION_NOT_QUEUED (_HRESULT_TYPEDEF_(0x80110600L))
value COMQC_E_BAD_MESSAGE (_HRESULT_TYPEDEF_(0x80110604L))
value COMQC_E_NO_IPERSISTSTREAM (_HRESULT_TYPEDEF_(0x80110603L))
value COMQC_E_NO_QUEUEABLE_INTERFACES (_HRESULT_TYPEDEF_(0x80110601L))
value COMQC_E_QUEUING_SERVICE_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x80110602L))
value COMQC_E_UNAUTHENTICATED (_HRESULT_TYPEDEF_(0x80110605L))
value COMQC_E_UNTRUSTED_ENQUEUER (_HRESULT_TYPEDEF_(0x80110606L))
value COM_RIGHTS_ACTIVATE_LOCAL (8)
value COM_RIGHTS_ACTIVATE_REMOTE (16)
value COM_RIGHTS_EXECUTE (1)
value COM_RIGHTS_EXECUTE_LOCAL (2)
value COM_RIGHTS_EXECUTE_REMOTE (4)
value CONDITION_VARIABLE_INIT (RTL_CONDITION_VARIABLE_INIT)
value CONDITION_VARIABLE_LOCKMODE_SHARED (RTL_CONDITION_VARIABLE_LOCKMODE_SHARED)
value CONFIRMSAFETYACTION_LOADOBJECT (0x00000001)
value CONNDLG_CONN_POINT (0x00000002)
value CONNDLG_HIDE_BOX (0x00000008)
value CONNDLG_NOT_PERSIST (0x00000020)
value CONNDLG_PERSIST (0x00000010)
value CONNDLG_RO_PATH (0x00000001)
value CONNDLG_USE_MRU (0x00000004)
value CONNECT_CMD_SAVECRED (0x00001000)
value CONNECT_COMMANDLINE (0x00000800)
value CONNECT_CRED_RESET (0x00002000)
value CONNECT_CURRENT_MEDIA (0x00000200)
value CONNECT_DEFERRED (0x00000400)
value CONNECT_GLOBAL_MAPPING (0x00040000)
value CONNECT_INTERACTIVE (0x00000008)
value CONNECT_LOCALDRIVE (0x00000100)
value CONNECT_NEED_DRIVE (0x00000020)
value CONNECT_PROMPT (0x00000010)
value CONNECT_REDIRECT (0x00000080)
value CONNECT_REFCOUNT (0x00000040)
value CONNECT_REQUIRE_INTEGRITY (0x00004000)
value CONNECT_REQUIRE_PRIVACY (0x00008000)
value CONNECT_RESERVED (0xFF000000)
value CONNECT_TEMPORARY (0x00000004)
value CONNECT_UPDATE_PROFILE (0x00000001)
value CONNECT_UPDATE_RECENT (0x00000002)
value CONNECT_WRITE_THROUGH_SEMANTICS (0x00010000)
value CONSOLE_CARET_SELECTION (0x0001)
value CONSOLE_CARET_VISIBLE (0x0002)
value CONSOLE_FULLSCREEN (1)
value CONSOLE_FULLSCREEN_HARDWARE (2)
value CONSOLE_FULLSCREEN_MODE (1)
value CONSOLE_MOUSE_DOWN (0x0008)
value CONSOLE_MOUSE_SELECTION (0x0004)
value CONSOLE_NO_SELECTION (0x0000)
value CONSOLE_SELECTION_IN_PROGRESS (0x0001)
value CONSOLE_SELECTION_NOT_EMPTY (0x0002)
value CONSOLE_TEXTMODE_BUFFER (1)
value CONSOLE_WINDOWED_MODE (2)
value CONTACTVISUALIZATION_OFF (0x0000)
value CONTACTVISUALIZATION_ON (0x0001)
value CONTACTVISUALIZATION_PRESENTATIONMODE (0x0002)
value CONTAINER_INHERIT_ACE ((0x2))
value CONTAINER_ROOT_INFO_FLAG_BIND_DO_NOT_MAP_NAME ((0x00000100))
value CONTAINER_ROOT_INFO_FLAG_BIND_EXCEPTION_ROOT ((0x00000080))
value CONTAINER_ROOT_INFO_FLAG_BIND_ROOT ((0x00000020))
value CONTAINER_ROOT_INFO_FLAG_BIND_TARGET_ROOT ((0x00000040))
value CONTAINER_ROOT_INFO_FLAG_LAYER_ROOT ((0x00000002))
value CONTAINER_ROOT_INFO_FLAG_SCRATCH_ROOT ((0x00000001))
value CONTAINER_ROOT_INFO_FLAG_UNION_LAYER_ROOT ((0x00000200))
value CONTAINER_ROOT_INFO_FLAG_VIRTUALIZATION_EXCEPTION_ROOT ((0x00000010))
value CONTAINER_ROOT_INFO_FLAG_VIRTUALIZATION_ROOT ((0x00000004))
value CONTAINER_ROOT_INFO_FLAG_VIRTUALIZATION_TARGET_ROOT ((0x00000008))
value CONTAINER_VOLUME_STATE_HOSTING_CONTAINER ((0x00000001))
value CONTEXT_ALL ((CONTEXT_CONTROL | CONTEXT_INTEGER | CONTEXT_SEGMENTS | CONTEXT_FLOATING_POINT | CONTEXT_DEBUG_REGISTERS))
value CONTEXT_CONTROL ((CONTEXT_AMD64 | 0x00000001L))
value CONTEXT_DEBUG_REGISTERS ((CONTEXT_AMD64 | 0x00000010L))
value CONTEXT_EXCEPTION_ACTIVE (0x08000000L)
value CONTEXT_EXCEPTION_REPORTING (0x80000000L)
value CONTEXT_EXCEPTION_REQUEST (0x40000000L)
value CONTEXT_E_ABORTED (_HRESULT_TYPEDEF_(0x8004E002L))
value CONTEXT_E_ABORTING (_HRESULT_TYPEDEF_(0x8004E003L))
value CONTEXT_E_FIRST (0x8004E000L)
value CONTEXT_E_LAST (0x8004E02FL)
value CONTEXT_E_NOCONTEXT (_HRESULT_TYPEDEF_(0x8004E004L))
value CONTEXT_E_NOJIT (_HRESULT_TYPEDEF_(0x8004E026L))
value CONTEXT_E_NOTRANSACTION (_HRESULT_TYPEDEF_(0x8004E027L))
value CONTEXT_E_OLDREF (_HRESULT_TYPEDEF_(0x8004E007L))
value CONTEXT_E_ROLENOTFOUND (_HRESULT_TYPEDEF_(0x8004E00CL))
value CONTEXT_E_SYNCH_TIMEOUT (_HRESULT_TYPEDEF_(0x8004E006L))
value CONTEXT_E_TMNOTAVAILABLE (_HRESULT_TYPEDEF_(0x8004E00FL))
value CONTEXT_E_WOULD_DEADLOCK (_HRESULT_TYPEDEF_(0x8004E005L))
value CONTEXT_FLOATING_POINT ((CONTEXT_AMD64 | 0x00000008L))
value CONTEXT_FULL ((CONTEXT_CONTROL | CONTEXT_INTEGER | CONTEXT_FLOATING_POINT))
value CONTEXT_INTEGER ((CONTEXT_AMD64 | 0x00000002L))
value CONTEXT_KERNEL_CET ((CONTEXT_AMD64 | 0x00000080L))
value CONTEXT_OID_CERTIFICATE (((LPCSTR)1))
value CONTEXT_OID_CRL (((LPCSTR)2))
value CONTEXT_OID_CTL (((LPCSTR)3))
value CONTEXT_OID_OCSP_RESP (((LPCSTR)6))
value CONTEXT_SEGMENTS ((CONTEXT_AMD64 | 0x00000004L))
value CONTEXT_SERVICE_ACTIVE (0x10000000L)
value CONTEXT_S_FIRST (0x0004E000L)
value CONTEXT_S_LAST (0x0004E02FL)
value CONTEXT_UNWOUND_TO_CALL (0x20000000)
value CONTEXT_XSTATE ((CONTEXT_AMD64 | 0x00000040L))
value CONTROL_C_EXIT (STATUS_CONTROL_C_EXIT)
value COPYFILE_SIS_FLAGS (0x0003)
value COPYFILE_SIS_LINK (0x0001)
value COPYFILE_SIS_REPLACE (0x0002)
value COPY_FILE_ALLOW_DECRYPTED_DESTINATION (0x00000008)
value COPY_FILE_COPY_SYMLINK (0x00000800)
value COPY_FILE_DIRECTORY (0x00000080)
value COPY_FILE_DISABLE_PRE_ALLOCATION (0x04000000)
value COPY_FILE_DONT_REQUEST_DEST_WRITE_DAC (0x02000000)
value COPY_FILE_ENABLE_LOW_FREE_SPACE_MODE (0x08000000)
value COPY_FILE_ENABLE_SPARSE_COPY (0x20000000)
value COPY_FILE_FAIL_IF_EXISTS (0x00000001)
value COPY_FILE_IGNORE_EDP_BLOCK (0x00400000)
value COPY_FILE_IGNORE_SOURCE_ENCRYPTION (0x00800000)
value COPY_FILE_NO_BUFFERING (0x00001000)
value COPY_FILE_NO_OFFLOAD (0x00040000)
value COPY_FILE_OPEN_AND_COPY_REPARSE_POINT (0x00200000)
value COPY_FILE_OPEN_SOURCE_FOR_WRITE (0x00000004)
value COPY_FILE_REQUEST_COMPRESSED_TRAFFIC (0x10000000)
value COPY_FILE_REQUEST_SECURITY_PRIVILEGES (0x00002000)
value COPY_FILE_RESTARTABLE (0x00000002)
value COPY_FILE_RESUME_FROM_PAUSE (0x00004000)
value COPY_FILE_SKIP_ALTERNATE_STREAMS (0x00008000)
value CORE_PARKING_POLICY_CHANGE_IDEAL (0)
value CORE_PARKING_POLICY_CHANGE_MAX (CORE_PARKING_POLICY_CHANGE_MULTISTEP)
value CORE_PARKING_POLICY_CHANGE_MULTISTEP (3)
value CORE_PARKING_POLICY_CHANGE_ROCKET (2)
value CORE_PARKING_POLICY_CHANGE_SINGLE (1)
value CO_E_ACCESSCHECKFAILED (_HRESULT_TYPEDEF_(0x8001012AL))
value CO_E_ACESINWRONGORDER (_HRESULT_TYPEDEF_(0x8001013AL))
value CO_E_ACNOTINITIALIZED (_HRESULT_TYPEDEF_(0x8001013FL))
value CO_E_ACTIVATIONFAILED (_HRESULT_TYPEDEF_(0x8004E021L))
value CO_E_ACTIVATIONFAILED_CATALOGERROR (_HRESULT_TYPEDEF_(0x8004E023L))
value CO_E_ACTIVATIONFAILED_EVENTLOGGED (_HRESULT_TYPEDEF_(0x8004E022L))
value CO_E_ACTIVATIONFAILED_TIMEOUT (_HRESULT_TYPEDEF_(0x8004E024L))
value CO_E_ALREADYINITIALIZED (_HRESULT_TYPEDEF_(0x800401F1L))
value CO_E_APPDIDNTREG (_HRESULT_TYPEDEF_(0x800401FEL))
value CO_E_APPNOTFOUND (_HRESULT_TYPEDEF_(0x800401F5L))
value CO_E_APPSINGLEUSE (_HRESULT_TYPEDEF_(0x800401F6L))
value CO_E_ASYNC_WORK_REJECTED (_HRESULT_TYPEDEF_(0x80004029L))
value CO_E_ATTEMPT_TO_CREATE_OUTSIDE_CLIENT_CONTEXT (_HRESULT_TYPEDEF_(0x80004024L))
value CO_E_BAD_PATH (_HRESULT_TYPEDEF_(0x80080004L))
value CO_E_BAD_SERVER_NAME (_HRESULT_TYPEDEF_(0x80004014L))
value CO_E_CALL_OUT_OF_TX_SCOPE_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x8004E030L))
value CO_E_CANCEL_DISABLED (_HRESULT_TYPEDEF_(0x80010140L))
value CO_E_CANTDETERMINECLASS (_HRESULT_TYPEDEF_(0x800401F2L))
value CO_E_CANT_REMOTE (_HRESULT_TYPEDEF_(0x80004013L))
value CO_E_CLASSSTRING (_HRESULT_TYPEDEF_(0x800401F3L))
value CO_E_CLASS_CREATE_FAILED (_HRESULT_TYPEDEF_(0x80080001L))
value CO_E_CLASS_DISABLED (_HRESULT_TYPEDEF_(0x80004027L))
value CO_E_CLRNOTAVAILABLE (_HRESULT_TYPEDEF_(0x80004028L))
value CO_E_CLSREG_INCONSISTENT (_HRESULT_TYPEDEF_(0x8000401FL))
value CO_E_CONVERSIONFAILED (_HRESULT_TYPEDEF_(0x8001012EL))
value CO_E_CREATEPROCESS_FAILURE (_HRESULT_TYPEDEF_(0x80004018L))
value CO_E_DBERROR (_HRESULT_TYPEDEF_(0x8004E02BL))
value CO_E_DECODEFAILED (_HRESULT_TYPEDEF_(0x8001013DL))
value CO_E_DLLNOTFOUND (_HRESULT_TYPEDEF_(0x800401F8L))
value CO_E_ELEVATION_DISABLED (_HRESULT_TYPEDEF_(0x80080017L))
value CO_E_ERRORINAPP (_HRESULT_TYPEDEF_(0x800401F7L))
value CO_E_ERRORINDLL (_HRESULT_TYPEDEF_(0x800401F9L))
value CO_E_EXCEEDSYSACLLIMIT (_HRESULT_TYPEDEF_(0x80010139L))
value CO_E_EXIT_TRANSACTION_SCOPE_NOT_CALLED (_HRESULT_TYPEDEF_(0x8004E031L))
value CO_E_FAILEDTOCLOSEHANDLE (_HRESULT_TYPEDEF_(0x80010138L))
value CO_E_FAILEDTOCREATEFILE (_HRESULT_TYPEDEF_(0x80010137L))
value CO_E_FAILEDTOGENUUID (_HRESULT_TYPEDEF_(0x80010136L))
value CO_E_FAILEDTOGETSECCTX (_HRESULT_TYPEDEF_(0x80010124L))
value CO_E_FAILEDTOGETTOKENINFO (_HRESULT_TYPEDEF_(0x80010126L))
value CO_E_FAILEDTOGETWINDIR (_HRESULT_TYPEDEF_(0x80010134L))
value CO_E_FAILEDTOIMPERSONATE (_HRESULT_TYPEDEF_(0x80010123L))
value CO_E_FAILEDTOOPENPROCESSTOKEN (_HRESULT_TYPEDEF_(0x8001013CL))
value CO_E_FAILEDTOOPENTHREADTOKEN (_HRESULT_TYPEDEF_(0x80010125L))
value CO_E_FAILEDTOQUERYCLIENTBLANKET (_HRESULT_TYPEDEF_(0x80010128L))
value CO_E_FAILEDTOSETDACL (_HRESULT_TYPEDEF_(0x80010129L))
value CO_E_FIRST (0x800401F0L)
value CO_E_IIDREG_INCONSISTENT (_HRESULT_TYPEDEF_(0x80004020L))
value CO_E_IIDSTRING (_HRESULT_TYPEDEF_(0x800401F4L))
value CO_E_INCOMPATIBLESTREAMVERSION (_HRESULT_TYPEDEF_(0x8001013BL))
value CO_E_INITIALIZATIONFAILED (_HRESULT_TYPEDEF_(0x8004E025L))
value CO_E_INIT_CLASS_CACHE (_HRESULT_TYPEDEF_(0x80004009L))
value CO_E_INIT_MEMORY_ALLOCATOR (_HRESULT_TYPEDEF_(0x80004008L))
value CO_E_INIT_ONLY_SINGLE_THREADED (_HRESULT_TYPEDEF_(0x80004012L))
value CO_E_INIT_RPC_CHANNEL (_HRESULT_TYPEDEF_(0x8000400AL))
value CO_E_INIT_SCM_EXEC_FAILURE (_HRESULT_TYPEDEF_(0x80004011L))
value CO_E_INIT_SCM_FILE_MAPPING_EXISTS (_HRESULT_TYPEDEF_(0x8000400FL))
value CO_E_INIT_SCM_MAP_VIEW_OF_FILE (_HRESULT_TYPEDEF_(0x80004010L))
value CO_E_INIT_SCM_MUTEX_EXISTS (_HRESULT_TYPEDEF_(0x8000400EL))
value CO_E_INIT_SHARED_ALLOCATOR (_HRESULT_TYPEDEF_(0x80004007L))
value CO_E_INIT_TLS (_HRESULT_TYPEDEF_(0x80004006L))
value CO_E_INIT_TLS_CHANNEL_CONTROL (_HRESULT_TYPEDEF_(0x8000400CL))
value CO_E_INIT_TLS_SET_CHANNEL_CONTROL (_HRESULT_TYPEDEF_(0x8000400BL))
value CO_E_INIT_UNACCEPTED_USER_ALLOCATOR (_HRESULT_TYPEDEF_(0x8000400DL))
value CO_E_INVALIDSID (_HRESULT_TYPEDEF_(0x8001012DL))
value CO_E_ISOLEVELMISMATCH (_HRESULT_TYPEDEF_(0x8004E02FL))
value CO_E_LAST (0x800401FFL)
value CO_E_LAUNCH_PERMSSION_DENIED (_HRESULT_TYPEDEF_(0x8000401BL))
value CO_E_LOOKUPACCNAMEFAILED (_HRESULT_TYPEDEF_(0x80010132L))
value CO_E_LOOKUPACCSIDFAILED (_HRESULT_TYPEDEF_(0x80010130L))
value CO_E_MALFORMED_SPN (_HRESULT_TYPEDEF_(0x80004033L))
value CO_E_MISSING_DISPLAYNAME (_HRESULT_TYPEDEF_(0x80080015L))
value CO_E_MSI_ERROR (_HRESULT_TYPEDEF_(0x80004023L))
value CO_E_NETACCESSAPIFAILED (_HRESULT_TYPEDEF_(0x8001012BL))
value CO_E_NOCOOKIES (_HRESULT_TYPEDEF_(0x8004E02AL))
value CO_E_NOIISINTRINSICS (_HRESULT_TYPEDEF_(0x8004E029L))
value CO_E_NOMATCHINGNAMEFOUND (_HRESULT_TYPEDEF_(0x80010131L))
value CO_E_NOMATCHINGSIDFOUND (_HRESULT_TYPEDEF_(0x8001012FL))
value CO_E_NOSYNCHRONIZATION (_HRESULT_TYPEDEF_(0x8004E02EL))
value CO_E_NOTCONSTRUCTED (_HRESULT_TYPEDEF_(0x8004E02DL))
value CO_E_NOTINITIALIZED (_HRESULT_TYPEDEF_(0x800401F0L))
value CO_E_NOTPOOLED (_HRESULT_TYPEDEF_(0x8004E02CL))
value CO_E_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80004021L))
value CO_E_NO_SECCTX_IN_ACTIVATE (_HRESULT_TYPEDEF_(0x8000402BL))
value CO_E_OBJISREG (_HRESULT_TYPEDEF_(0x800401FCL))
value CO_E_OBJNOTCONNECTED (_HRESULT_TYPEDEF_(0x800401FDL))
value CO_E_OBJNOTREG (_HRESULT_TYPEDEF_(0x800401FBL))
value CO_E_OBJSRV_RPC_FAILURE (_HRESULT_TYPEDEF_(0x80080006L))
value CO_E_PATHTOOLONG (_HRESULT_TYPEDEF_(0x80010135L))
value CO_E_PREMATURE_STUB_RUNDOWN (_HRESULT_TYPEDEF_(0x80004035L))
value CO_E_RELEASED (_HRESULT_TYPEDEF_(0x800401FFL))
value CO_E_RELOAD_DLL (_HRESULT_TYPEDEF_(0x80004022L))
value CO_E_REMOTE_COMMUNICATION_FAILURE (_HRESULT_TYPEDEF_(0x8000401DL))
value CO_E_RUNAS_CREATEPROCESS_FAILURE (_HRESULT_TYPEDEF_(0x80004019L))
value CO_E_RUNAS_LOGON_FAILURE (_HRESULT_TYPEDEF_(0x8000401AL))
value CO_E_RUNAS_SYNTAX (_HRESULT_TYPEDEF_(0x80004017L))
value CO_E_RUNAS_VALUE_MUST_BE_AAA (_HRESULT_TYPEDEF_(0x80080016L))
value CO_E_SCM_ERROR (_HRESULT_TYPEDEF_(0x80080002L))
value CO_E_SCM_RPC_FAILURE (_HRESULT_TYPEDEF_(0x80080003L))
value CO_E_SERVER_EXEC_FAILURE (_HRESULT_TYPEDEF_(0x80080005L))
value CO_E_SERVER_INIT_TIMEOUT (_HRESULT_TYPEDEF_(0x8000402AL))
value CO_E_SERVER_NOT_PAUSED (_HRESULT_TYPEDEF_(0x80004026L))
value CO_E_SERVER_PAUSED (_HRESULT_TYPEDEF_(0x80004025L))
value CO_E_SERVER_START_TIMEOUT (_HRESULT_TYPEDEF_(0x8000401EL))
value CO_E_SERVER_STOPPING (_HRESULT_TYPEDEF_(0x80080008L))
value CO_E_SETSERLHNDLFAILED (_HRESULT_TYPEDEF_(0x80010133L))
value CO_E_START_SERVICE_FAILURE (_HRESULT_TYPEDEF_(0x8000401CL))
value CO_E_SXS_CONFIG (_HRESULT_TYPEDEF_(0x80004032L))
value CO_E_THREADINGMODEL_CHANGED (_HRESULT_TYPEDEF_(0x8004E028L))
value CO_E_THREADPOOL_CONFIG (_HRESULT_TYPEDEF_(0x80004031L))
value CO_E_TRACKER_CONFIG (_HRESULT_TYPEDEF_(0x80004030L))
value CO_E_TRUSTEEDOESNTMATCHCLIENT (_HRESULT_TYPEDEF_(0x80010127L))
value CO_E_UNREVOKED_REGISTRATION_ON_APARTMENT_SHUTDOWN (_HRESULT_TYPEDEF_(0x80004034L))
value CO_E_WRONGOSFORAPP (_HRESULT_TYPEDEF_(0x800401FAL))
value CO_E_WRONGTRUSTEENAMESYNTAX (_HRESULT_TYPEDEF_(0x8001012CL))
value CO_E_WRONG_SERVER_IDENTITY (_HRESULT_TYPEDEF_(0x80004015L))
value CO_S_FIRST (0x000401F0L)
value CO_S_LAST (0x000401FFL)
value CO_S_MACHINENAMENOTFOUND (_HRESULT_TYPEDEF_(0x00080013L))
value CO_S_NOTALLINTERFACES (_HRESULT_TYPEDEF_(0x00080012L))
value CPS_CANCEL (0x0004)
value CPS_COMPLETE (0x0001)
value CPS_CONVERT (0x0002)
value CPS_REVERT (0x0003)
value CP_ACP (0)
value CP_INSTALLED (0x00000001)
value CP_MACCP (2)
value CP_NONE (0)
value CP_OEMCP (1)
value CP_RECTANGLE (1)
value CP_REGION (2)
value CP_SUPPORTED (0x00000002)
value CP_SYMBOL (42)
value CP_THREAD_ACP (3)
value CP_WINANSI (1004)
value CP_WINNEUTRAL (CP_WINANSI)
value CP_WINUNICODE (1200)
value CREATECOLORSPACE_EMBEDED (0x00000001)
value CREATEPROCESS_MANIFEST_RESOURCE_ID (MAKEINTRESOURCE( 1))
value CREATE_ALWAYS (2)
value CREATE_BOUNDARY_DESCRIPTOR_ADD_APPCONTAINER_SID (0x1)
value CREATE_BREAKAWAY_FROM_JOB (0x01000000)
value CREATE_DEFAULT_ERROR_MODE (0x04000000)
value CREATE_EVENT_INITIAL_SET (0x00000002)
value CREATE_EVENT_MANUAL_RESET (0x00000001)
value CREATE_FORCEDOS (0x00002000)
value CREATE_FOR_DIR ((2))
value CREATE_FOR_IMPORT ((1))
value CREATE_IGNORE_SYSTEM_DEFAULT (0x80000000)
value CREATE_MUTEX_INITIAL_OWNER (0x00000001)
value CREATE_NEW (1)
value CREATE_NEW_CONSOLE (0x00000010)
value CREATE_NEW_PROCESS_GROUP (0x00000200)
value CREATE_NO_WINDOW (0x08000000)
value CREATE_PRESERVE_CODE_AUTHZ_LEVEL (0x02000000)
value CREATE_PROCESS_DEBUG_EVENT (3)
value CREATE_PROTECTED_PROCESS (0x00040000)
value CREATE_SECURE_PROCESS (0x00400000)
value CREATE_SEPARATE_WOW_VDM (0x00000800)
value CREATE_SHARED_WOW_VDM (0x00001000)
value CREATE_SUSPENDED (0x00000004)
value CREATE_THREAD_DEBUG_EVENT (2)
value CREATE_UNICODE_ENVIRONMENT (0x00000400)
value CREATE_WAITABLE_TIMER_HIGH_RESOLUTION (0x00000002)
value CREATE_WAITABLE_TIMER_MANUAL_RESET (0x00000001)
value CREDENTIAL_OID_PASSWORD_CREDENTIALS (CREDENTIAL_OID_PASSWORD_CREDENTIALS_A)
value CREDENTIAL_OID_PASSWORD_CREDENTIALS_A (((LPCSTR)1))
value CREDENTIAL_OID_PASSWORD_CREDENTIALS_W (((LPCSTR)2))
value CRITICAL_ACE_FLAG ((0x20))
value CRITICAL_SECTION_NO_DEBUG_INFO (RTL_CRITICAL_SECTION_FLAG_NO_DEBUG_INFO)
value CRL_DIST_POINT_ERR_CRL_ISSUER_BIT (0x80000000L)
value CRL_DIST_POINT_ERR_INDEX_MASK (0x7F)
value CRL_DIST_POINT_ERR_INDEX_SHIFT (24)
value CRL_DIST_POINT_FULL_NAME (1)
value CRL_DIST_POINT_ISSUER_RDN_NAME (2)
value CRL_DIST_POINT_NO_NAME (0)
value CRL_FIND_ANY (0)
value CRL_FIND_EXISTING (2)
value CRL_FIND_ISSUED_BY (1)
value CRL_FIND_ISSUED_BY_AKI_FLAG (0x1)
value CRL_FIND_ISSUED_BY_BASE_FLAG (0x8)
value CRL_FIND_ISSUED_BY_DELTA_FLAG (0x4)
value CRL_FIND_ISSUED_BY_SIGNATURE_FLAG (0x2)
value CRL_FIND_ISSUED_FOR (3)
value CRL_FIND_ISSUED_FOR_SET_STRONG_PROPERTIES_FLAG (0x10)
value CRL_REASON_AA_COMPROMISE (10)
value CRL_REASON_AA_COMPROMISE_FLAG (0x80)
value CRL_REASON_AFFILIATION_CHANGED (3)
value CRL_REASON_AFFILIATION_CHANGED_FLAG (0x10)
value CRL_REASON_CA_COMPROMISE (2)
value CRL_REASON_CA_COMPROMISE_FLAG (0x20)
value CRL_REASON_CERTIFICATE_HOLD (6)
value CRL_REASON_CERTIFICATE_HOLD_FLAG (0x02)
value CRL_REASON_CESSATION_OF_OPERATION (5)
value CRL_REASON_CESSATION_OF_OPERATION_FLAG (0x04)
value CRL_REASON_KEY_COMPROMISE (1)
value CRL_REASON_KEY_COMPROMISE_FLAG (0x40)
value CRL_REASON_PRIVILEGE_WITHDRAWN (9)
value CRL_REASON_PRIVILEGE_WITHDRAWN_FLAG (0x01)
value CRL_REASON_REMOVE_FROM_CRL (8)
value CRL_REASON_SUPERSEDED (4)
value CRL_REASON_SUPERSEDED_FLAG (0x08)
value CRL_REASON_UNSPECIFIED (0)
value CRL_REASON_UNUSED_FLAG (0x80)
value CRM_PROTOCOL_DYNAMIC_MARSHAL_INFO (0x00000002)
value CRM_PROTOCOL_EXPLICIT_MARSHAL_ONLY (0x00000001)
value CRM_PROTOCOL_MAXIMUM_OPTION (0x00000003)
value CROSS_CERT_DIST_POINT_ERR_INDEX_MASK (0xFF)
value CROSS_CERT_DIST_POINT_ERR_INDEX_SHIFT (24)
value CRYPTNET_CACHED_OCSP_SWITCH_TO_CRL_COUNT_DEFAULT (50)
value CRYPTNET_CRL_BEFORE_OCSP_ENABLE (0xFFFFFFFF)
value CRYPTNET_MAX_CACHED_OCSP_PER_CRL_COUNT_DEFAULT (500)
value CRYPTNET_OCSP_AFTER_CRL_DISABLE (0xFFFFFFFF)
value CRYPTNET_PRE_FETCH_AFTER_PUBLISH_PRE_FETCH_DIVISOR_DEFAULT (10)
value CRYPTNET_PRE_FETCH_BEFORE_NEXT_UPDATE_PRE_FETCH_DIVISOR_DEFAULT (20)
value CRYPTNET_PRE_FETCH_SCAN_AFTER_TRIGGER_DELAY_SECONDS_DEFAULT (60)
value CRYPTNET_PRE_FETCH_TRIGGER_DISABLE (0xFFFFFFFF)
value CRYPTNET_PRE_FETCH_VALIDITY_PERIOD_AFTER_NEXT_UPDATE_PRE_FETCH_DIVISOR_DEFAULT (10)
value CRYPTNET_URL_CACHE_DEFAULT_FLUSH (0)
value CRYPTNET_URL_CACHE_DISABLE_FLUSH (0xFFFFFFFF)
value CRYPTNET_URL_CACHE_PRE_FETCH_AUTOROOT_CAB (5)
value CRYPTNET_URL_CACHE_PRE_FETCH_BLOB (1)
value CRYPTNET_URL_CACHE_PRE_FETCH_CRL (2)
value CRYPTNET_URL_CACHE_PRE_FETCH_DISALLOWED_CERT_CAB (6)
value CRYPTNET_URL_CACHE_PRE_FETCH_NONE (0)
value CRYPTNET_URL_CACHE_PRE_FETCH_OCSP (3)
value CRYPTNET_URL_CACHE_PRE_FETCH_PIN_RULES_CAB (7)
value CRYPTNET_URL_CACHE_RESPONSE_HTTP (1)
value CRYPTNET_URL_CACHE_RESPONSE_NONE (0)
value CRYPTNET_URL_CACHE_RESPONSE_VALIDATED (0x8000)
value CRYPTPROTECTMEMORY_BLOCK_SIZE (16)
value CRYPTPROTECTMEMORY_CROSS_PROCESS (0x01)
value CRYPTPROTECTMEMORY_SAME_LOGON (0x02)
value CRYPTPROTECTMEMORY_SAME_PROCESS (0x00)
value CRYPTPROTECT_AUDIT (0x10)
value CRYPTPROTECT_CRED_REGENERATE (0x80)
value CRYPTPROTECT_CRED_SYNC (0x8)
value CRYPTPROTECT_FIRST_RESERVED_FLAGVAL (0x0FFFFFFF)
value CRYPTPROTECT_LAST_RESERVED_FLAGVAL (0xFFFFFFFF)
value CRYPTPROTECT_LOCAL_MACHINE (0x4)
value CRYPTPROTECT_NO_RECOVERY (0x20)
value CRYPTPROTECT_PROMPT_ON_PROTECT (0x2)
value CRYPTPROTECT_PROMPT_ON_UNPROTECT (0x1)
value CRYPTPROTECT_PROMPT_REQUIRE_STRONG (0x10)
value CRYPTPROTECT_PROMPT_RESERVED (0x04)
value CRYPTPROTECT_PROMPT_STRONG (0x08)
value CRYPTPROTECT_UI_FORBIDDEN (0x1)
value CRYPTPROTECT_VERIFY_PROTECTION (0x40)
value CRYPT_ACCUMULATIVE_TIMEOUT (0x00000800)
value CRYPT_ACQUIRE_ALLOW_NCRYPT_KEY_FLAG (0x00010000)
value CRYPT_ACQUIRE_CACHE_FLAG (0x00000001)
value CRYPT_ACQUIRE_COMPARE_KEY_FLAG (0x00000004)
value CRYPT_ACQUIRE_NCRYPT_KEY_FLAGS_MASK (0x00070000)
value CRYPT_ACQUIRE_NO_HEALING (0x00000008)
value CRYPT_ACQUIRE_ONLY_NCRYPT_KEY_FLAG (0x00040000)
value CRYPT_ACQUIRE_PREFER_NCRYPT_KEY_FLAG (0x00020000)
value CRYPT_ACQUIRE_SILENT_FLAG (0x00000040)
value CRYPT_ACQUIRE_USE_PROV_INFO_FLAG (0x00000002)
value CRYPT_ACQUIRE_WINDOW_HANDLE_FLAG (0x00000080)
value CRYPT_AIA_RETRIEVAL (0x00080000)
value CRYPT_ALL_FUNCTIONS ((0x00000001))
value CRYPT_ALL_PROVIDERS ((0x00000002))
value CRYPT_ANY ((0x00000004))
value CRYPT_ARCHIVABLE (0x00004000)
value CRYPT_ARCHIVE (0x0100)
value CRYPT_ASN_ENCODING (0x00000001)
value CRYPT_ASYNC_RETRIEVAL (0x00000010)
value CRYPT_CACHE_ONLY_RETRIEVAL (0x00000002)
value CRYPT_CHECK_FRESHNESS_TIME_VALIDITY (0x00000400)
value CRYPT_CREATE_IV (0x00000200)
value CRYPT_CREATE_NEW_FLUSH_ENTRY (0x10000000)
value CRYPT_CREATE_SALT (0x00000004)
value CRYPT_DATA_KEY (0x00000800)
value CRYPT_DECODE_ALLOC_FLAG (0x8000)
value CRYPT_DECODE_ENABLE_PUNYCODE_FLAG (0x02000000)
value CRYPT_DECODE_NOCOPY_FLAG (0x1)
value CRYPT_DECODE_NO_SIGNATURE_BYTE_REVERSAL_FLAG (0x8)
value CRYPT_DECODE_SHARE_OID_STRING_FLAG (0x4)
value CRYPT_DECODE_TO_BE_SIGNED_FLAG (0x2)
value CRYPT_DECRYPT (0x0002)
value CRYPT_DECRYPT_RSA_NO_PADDING_CHECK (0x00000020)
value CRYPT_DEFAULT_CONTAINER_OPTIONAL (0x00000080)
value CRYPT_DEFAULT_CONTEXT_AUTO_RELEASE_FLAG (0x00000001)
value CRYPT_DEFAULT_CONTEXT_CERT_SIGN_OID (1)
value CRYPT_DEFAULT_CONTEXT_MULTI_CERT_SIGN_OID (2)
value CRYPT_DEFAULT_CONTEXT_PROCESS_FLAG (0x00000002)
value CRYPT_DELETEKEYSET (0x00000010)
value CRYPT_DELETE_DEFAULT (0x00000004)
value CRYPT_DELETE_KEYSET (CRYPT_DELETEKEYSET)
value CRYPT_DESTROYKEY (0x00000004)
value CRYPT_DOMAIN ((0x00000002))
value CRYPT_DONT_CACHE_RESULT (0x00000008)
value CRYPT_DONT_CHECK_TIME_VALIDITY (0x00000200)
value CRYPT_DONT_VERIFY_SIGNATURE (0x00000100)
value CRYPT_ECC_CMS_SHARED_INFO_SUPPPUBINFO_BYTE_LENGTH (4)
value CRYPT_ENABLE_FILE_RETRIEVAL (0x08000000)
value CRYPT_ENABLE_SSL_REVOCATION_RETRIEVAL (0x00800000)
value CRYPT_ENCODE_ALLOC_FLAG (0x8000)
value CRYPT_ENCODE_DECODE_NONE (0)
value CRYPT_ENCODE_ENABLE_PUNYCODE_FLAG (0x20000)
value CRYPT_ENCODE_NO_SIGNATURE_BYTE_REVERSAL_FLAG (0x8)
value CRYPT_ENCRYPT (0x0001)
value CRYPT_ENCRYPT_ALG_OID_GROUP_ID (2)
value CRYPT_ENHKEY_USAGE_OID_GROUP_ID (7)
value CRYPT_EXCLUSIVE ((0x00000001))
value CRYPT_EXPORT (0x0004)
value CRYPT_EXPORTABLE (0x00000001)
value CRYPT_EXPORT_KEY (0x0040)
value CRYPT_EXT_OR_ATTR_OID_GROUP_ID (6)
value CRYPT_E_ALREADY_DECRYPTED (_HRESULT_TYPEDEF_(0x80091009L))
value CRYPT_E_ATTRIBUTES_MISSING (_HRESULT_TYPEDEF_(0x8009100FL))
value CRYPT_E_AUTH_ATTR_MISSING (_HRESULT_TYPEDEF_(0x80091006L))
value CRYPT_E_BAD_ENCODE (_HRESULT_TYPEDEF_(0x80092002L))
value CRYPT_E_BAD_LEN (_HRESULT_TYPEDEF_(0x80092001L))
value CRYPT_E_BAD_MSG (_HRESULT_TYPEDEF_(0x8009200DL))
value CRYPT_E_CONTROL_TYPE (_HRESULT_TYPEDEF_(0x8009100CL))
value CRYPT_E_DELETED_PREV (_HRESULT_TYPEDEF_(0x80092008L))
value CRYPT_E_EXISTS (_HRESULT_TYPEDEF_(0x80092005L))
value CRYPT_E_FILERESIZED (_HRESULT_TYPEDEF_(0x80092025L))
value CRYPT_E_FILE_ERROR (_HRESULT_TYPEDEF_(0x80092003L))
value CRYPT_E_HASH_VALUE (_HRESULT_TYPEDEF_(0x80091007L))
value CRYPT_E_INVALID_INDEX (_HRESULT_TYPEDEF_(0x80091008L))
value CRYPT_E_INVALID_MSG_TYPE (_HRESULT_TYPEDEF_(0x80091004L))
value CRYPT_E_INVALID_NUMERIC_STRING (_HRESULT_TYPEDEF_(0x80092020L))
value CRYPT_E_INVALID_PRINTABLE_STRING (_HRESULT_TYPEDEF_(0x80092021L))
value CRYPT_E_ISSUER_SERIALNUMBER (_HRESULT_TYPEDEF_(0x8009100DL))
value CRYPT_E_MISSING_PUBKEY_PARA (_HRESULT_TYPEDEF_(0x8009202CL))
value CRYPT_E_MSG_ERROR (_HRESULT_TYPEDEF_(0x80091001L))
value CRYPT_E_NOT_CHAR_STRING (_HRESULT_TYPEDEF_(0x80092024L))
value CRYPT_E_NOT_DECRYPTED (_HRESULT_TYPEDEF_(0x8009100AL))
value CRYPT_E_NOT_FOUND (_HRESULT_TYPEDEF_(0x80092004L))
value CRYPT_E_NOT_IN_CTL (_HRESULT_TYPEDEF_(0x8009202AL))
value CRYPT_E_NOT_IN_REVOCATION_DATABASE (_HRESULT_TYPEDEF_(0x80092014L))
value CRYPT_E_NO_DECRYPT_CERT (_HRESULT_TYPEDEF_(0x8009200CL))
value CRYPT_E_NO_KEY_PROPERTY (_HRESULT_TYPEDEF_(0x8009200BL))
value CRYPT_E_NO_MATCH (_HRESULT_TYPEDEF_(0x80092009L))
value CRYPT_E_NO_PROVIDER (_HRESULT_TYPEDEF_(0x80092006L))
value CRYPT_E_NO_REVOCATION_CHECK (_HRESULT_TYPEDEF_(0x80092012L))
value CRYPT_E_NO_REVOCATION_DLL (_HRESULT_TYPEDEF_(0x80092011L))
value CRYPT_E_NO_SIGNER (_HRESULT_TYPEDEF_(0x8009200EL))
value CRYPT_E_NO_TRUSTED_SIGNER (_HRESULT_TYPEDEF_(0x8009202BL))
value CRYPT_E_NO_VERIFY_USAGE_CHECK (_HRESULT_TYPEDEF_(0x80092028L))
value CRYPT_E_NO_VERIFY_USAGE_DLL (_HRESULT_TYPEDEF_(0x80092027L))
value CRYPT_E_OBJECT_LOCATOR_OBJECT_NOT_FOUND (_HRESULT_TYPEDEF_(0x8009202DL))
value CRYPT_E_OID_FORMAT (_HRESULT_TYPEDEF_(0x80091003L))
value CRYPT_E_OSS_ERROR (_HRESULT_TYPEDEF_(0x80093000L))
value CRYPT_E_PENDING_CLOSE (_HRESULT_TYPEDEF_(0x8009200FL))
value CRYPT_E_RECIPIENT_NOT_FOUND (_HRESULT_TYPEDEF_(0x8009100BL))
value CRYPT_E_REVOCATION_OFFLINE (_HRESULT_TYPEDEF_(0x80092013L))
value CRYPT_E_REVOKED (_HRESULT_TYPEDEF_(0x80092010L))
value CRYPT_E_SECURITY_SETTINGS (_HRESULT_TYPEDEF_(0x80092026L))
value CRYPT_E_SELF_SIGNED (_HRESULT_TYPEDEF_(0x80092007L))
value CRYPT_E_SIGNER_NOT_FOUND (_HRESULT_TYPEDEF_(0x8009100EL))
value CRYPT_E_STREAM_INSUFFICIENT_DATA (_HRESULT_TYPEDEF_(0x80091011L))
value CRYPT_E_STREAM_MSG_NOT_READY (_HRESULT_TYPEDEF_(0x80091010L))
value CRYPT_E_UNEXPECTED_ENCODING (_HRESULT_TYPEDEF_(0x80091005L))
value CRYPT_E_UNEXPECTED_MSG_TYPE (_HRESULT_TYPEDEF_(0x8009200AL))
value CRYPT_E_UNKNOWN_ALGO (_HRESULT_TYPEDEF_(0x80091002L))
value CRYPT_E_VERIFY_USAGE_OFFLINE (_HRESULT_TYPEDEF_(0x80092029L))
value CRYPT_FAILED (FALSE)
value CRYPT_FASTSGC (0x0002)
value CRYPT_FIND_MACHINE_KEYSET_FLAG (0x00000002)
value CRYPT_FIND_SILENT_KEYSET_FLAG (0x00000040)
value CRYPT_FIND_USER_KEYSET_FLAG (0x00000001)
value CRYPT_FIRST (1)
value CRYPT_FIRST_ALG_OID_GROUP_ID (CRYPT_HASH_ALG_OID_GROUP_ID)
value CRYPT_FLAG_IPSEC (0x0010)
value CRYPT_FLAG_SIGNING (0x0020)
value CRYPT_FORCE_KEY_PROTECTION_HIGH (0x00008000)
value CRYPT_FORMAT_COMMA (0x1000)
value CRYPT_FORMAT_CRLF (CRYPT_FORMAT_RDN_CRLF)
value CRYPT_FORMAT_OID (0x0004)
value CRYPT_FORMAT_RDN_CRLF (0x0200)
value CRYPT_FORMAT_RDN_REVERSE (0x0800)
value CRYPT_FORMAT_RDN_SEMICOLON (0x0100)
value CRYPT_FORMAT_RDN_UNQUOTE (0x0400)
value CRYPT_FORMAT_SEMICOLON (CRYPT_FORMAT_RDN_SEMICOLON)
value CRYPT_FORMAT_SIMPLE (0x0001)
value CRYPT_FORMAT_STR_MULTI_LINE (0x0001)
value CRYPT_FORMAT_STR_NO_HEX (0x0010)
value CRYPT_GET_INSTALLED_OID_FUNC_FLAG (0x1)
value CRYPT_GET_URL_FROM_AUTH_ATTRIBUTE (0x00000008)
value CRYPT_GET_URL_FROM_EXTENSION (0x00000002)
value CRYPT_GET_URL_FROM_PROPERTY (0x00000001)
value CRYPT_GET_URL_FROM_UNAUTH_ATTRIBUTE (0x00000004)
value CRYPT_HASH_ALG_OID_GROUP_ID (1)
value CRYPT_HTTP_POST_RETRIEVAL (0x00100000)
value CRYPT_IMPL_HARDWARE (1)
value CRYPT_IMPL_MIXED (3)
value CRYPT_IMPL_REMOVABLE (8)
value CRYPT_IMPL_SOFTWARE (2)
value CRYPT_IMPL_UNKNOWN (4)
value CRYPT_IMPORT_KEY (0x0080)
value CRYPT_INITIATOR (0x00000040)
value CRYPT_INSTALL_OID_FUNC_BEFORE_FLAG (1)
value CRYPT_INSTALL_OID_INFO_BEFORE_FLAG (1)
value CRYPT_IPSEC_HMAC_KEY (0x00000100)
value CRYPT_I_NEW_PROTECTION_REQUIRED (_HRESULT_TYPEDEF_(0x00091012L))
value CRYPT_KDF_OID_GROUP_ID (10)
value CRYPT_KEEP_TIME_VALID (0x00000080)
value CRYPT_KEK (0x00000400)
value CRYPT_KEYID_ALLOC_FLAG (0x00008000)
value CRYPT_KEYID_DELETE_FLAG (0x00000010)
value CRYPT_KEYID_MACHINE_FLAG (0x00000020)
value CRYPT_KEYID_SET_NEW_FLAG (0x00002000)
value CRYPT_KM ((0x00000002))
value CRYPT_LAST_ALG_OID_GROUP_ID (CRYPT_SIGN_ALG_OID_GROUP_ID)
value CRYPT_LAST_OID_GROUP_ID (10)
value CRYPT_LDAP_AREC_EXCLUSIVE_RETRIEVAL (0x00040000)
value CRYPT_LDAP_INSERT_ENTRY_ATTRIBUTE (0x00008000)
value CRYPT_LDAP_SCOPE_BASE_ONLY_RETRIEVAL (0x00002000)
value CRYPT_LDAP_SIGN_RETRIEVAL (0x00010000)
value CRYPT_LITTLE_ENDIAN (0x00000001)
value CRYPT_LOCAL ((0x00000001))
value CRYPT_LOCALIZED_NAME_ENCODING_TYPE (0)
value CRYPT_MAC (0x0020)
value CRYPT_MACHINE_DEFAULT (0x00000001)
value CRYPT_MACHINE_KEYSET (0x00000020)
value CRYPT_MATCH_ANY_ENCODING_TYPE (0xFFFFFFFF)
value CRYPT_MESSAGE_BARE_CONTENT_OUT_FLAG (0x00000001)
value CRYPT_MESSAGE_ENCAPSULATED_CONTENT_OUT_FLAG (0x00000002)
value CRYPT_MESSAGE_KEYID_RECIPIENT_FLAG (0x4)
value CRYPT_MESSAGE_KEYID_SIGNER_FLAG (0x00000004)
value CRYPT_MESSAGE_SILENT_KEYSET_FLAG (0x00000040)
value CRYPT_MIN_DEPENDENCIES ((0x00000001))
value CRYPT_MM ((0x00000003))
value CRYPT_MODE_CBC (1)
value CRYPT_MODE_CBCI (6)
value CRYPT_MODE_CBCOFM (9)
value CRYPT_MODE_CBCOFMI (10)
value CRYPT_MODE_CFB (4)
value CRYPT_MODE_CFBP (7)
value CRYPT_MODE_CTS (5)
value CRYPT_MODE_ECB (2)
value CRYPT_MODE_OFB (3)
value CRYPT_MODE_OFBP (8)
value CRYPT_NDR_ENCODING (0x00000002)
value CRYPT_NEWKEYSET (0x00000008)
value CRYPT_NEXT (2)
value CRYPT_NOHASHOID (0x00000001)
value CRYPT_NOT_MODIFIED_RETRIEVAL (0x00400000)
value CRYPT_NO_AUTH_RETRIEVAL (0x00020000)
value CRYPT_NO_OCSP_FAILOVER_TO_CRL_RETRIEVAL (0x02000000)
value CRYPT_NO_SALT (0x00000010)
value CRYPT_OAEP (0x00000040)
value CRYPT_OBJECT_LOCATOR_FIRST_RESERVED_USER_NAME_TYPE (33)
value CRYPT_OBJECT_LOCATOR_LAST_RESERVED_NAME_TYPE (32)
value CRYPT_OBJECT_LOCATOR_LAST_RESERVED_USER_NAME_TYPE (0x0000FFFF)
value CRYPT_OBJECT_LOCATOR_RELEASE_DLL_UNLOAD (4)
value CRYPT_OBJECT_LOCATOR_RELEASE_PROCESS_EXIT (3)
value CRYPT_OBJECT_LOCATOR_RELEASE_SERVICE_STOP (2)
value CRYPT_OBJECT_LOCATOR_RELEASE_SYSTEM_SHUTDOWN (1)
value CRYPT_OBJECT_LOCATOR_SPN_NAME_TYPE (1)
value CRYPT_OCSP_ONLY_RETRIEVAL (0x01000000)
value CRYPT_OFFLINE_CHECK_RETRIEVAL (0x00004000)
value CRYPT_OID_DISABLE_SEARCH_DS_FLAG (0x80000000)
value CRYPT_OID_INFO_ALGID_KEY (3)
value CRYPT_OID_INFO_CNG_ALGID_KEY (5)
value CRYPT_OID_INFO_CNG_SIGN_KEY (6)
value CRYPT_OID_INFO_NAME_KEY (2)
value CRYPT_OID_INFO_OID_GROUP_BIT_LEN_MASK (0x0FFF0000)
value CRYPT_OID_INFO_OID_GROUP_BIT_LEN_SHIFT (16)
value CRYPT_OID_INFO_OID_KEY (1)
value CRYPT_OID_INFO_OID_KEY_FLAGS_MASK (0xFFFF0000)
value CRYPT_OID_INFO_PUBKEY_ENCRYPT_KEY_FLAG (0x40000000)
value CRYPT_OID_INFO_PUBKEY_SIGN_KEY_FLAG (0x80000000)
value CRYPT_OID_INFO_SIGN_KEY (4)
value CRYPT_OID_INHIBIT_SIGNATURE_FORMAT_FLAG (0x00000001)
value CRYPT_OID_NO_NULL_ALGORITHM_PARA_FLAG (0x00000004)
value CRYPT_OID_PUBKEY_ENCRYPT_ONLY_FLAG (0x40000000)
value CRYPT_OID_PUBKEY_SIGN_ONLY_FLAG (0x80000000)
value CRYPT_OID_USE_CURVE_NAME_FOR_ENCODE_FLAG (0x20000000)
value CRYPT_OID_USE_CURVE_PARAMETERS_FOR_ENCODE_FLAG (0x10000000)
value CRYPT_ONLINE (0x00000080)
value CRYPT_OVERRIDE ((0x00010000))
value CRYPT_OVERWRITE ((0x00000001))
value CRYPT_OWF_REPL_LM_HASH (0x00000001)
value CRYPT_PARAM_ASYNC_RETRIEVAL_COMPLETION (((LPCSTR)1))
value CRYPT_PARAM_CANCEL_ASYNC_RETRIEVAL (((LPCSTR)2))
value CRYPT_POLICY_OID_GROUP_ID (8)
value CRYPT_PREGEN (0x00000040)
value CRYPT_PRIORITY_BOTTOM ((0xFFFFFFFF))
value CRYPT_PRIORITY_TOP ((0x00000000))
value CRYPT_PROCESS_ISOLATE ((0x00010000))
value CRYPT_PROXY_CACHE_RETRIEVAL (0x00200000)
value CRYPT_PSTORE (0x00000002)
value CRYPT_PUBKEY_ALG_OID_GROUP_ID (3)
value CRYPT_RANDOM_QUERY_STRING_RETRIEVAL (0x04000000)
value CRYPT_RDN_ATTR_OID_GROUP_ID (5)
value CRYPT_READ (0x0008)
value CRYPT_RECIPIENT (0x00000010)
value CRYPT_REGISTER_FIRST_INDEX (0)
value CRYPT_REGISTER_LAST_INDEX (0xFFFFFFFF)
value CRYPT_RETRIEVE_MAX_ERROR_CONTENT_LENGTH (0x1000)
value CRYPT_RETRIEVE_MULTIPLE_OBJECTS (0x00000001)
value CRYPT_SECRETDIGEST (0x00000001)
value CRYPT_SEC_DESCR (0x00000001)
value CRYPT_SERVER (0x00000400)
value CRYPT_SF (0x00000100)
value CRYPT_SGC (0x0001)
value CRYPT_SGCKEY (0x00002000)
value CRYPT_SGC_ENUM (4)
value CRYPT_SIGN_ALG_OID_GROUP_ID (4)
value CRYPT_SILENT (0x00000040)
value CRYPT_SORTED_CTL_ENCODE_HASHED_SUBJECT_IDENTIFIER_FLAG (0x10000)
value CRYPT_STICKY_CACHE_RETRIEVAL (0x00001000)
value CRYPT_STRING_ANY (0x00000007)
value CRYPT_STRING_BINARY (0x00000002)
value CRYPT_STRING_ENCODEMASK (0x000000ff)
value CRYPT_STRING_HASHDATA (0x10000000)
value CRYPT_STRING_HEX (0x00000004)
value CRYPT_STRING_HEXADDR (0x0000000a)
value CRYPT_STRING_HEXASCII (0x00000005)
value CRYPT_STRING_HEXASCIIADDR (0x0000000b)
value CRYPT_STRING_HEXRAW (0x0000000c)
value CRYPT_STRING_HEX_ANY (0x00000008)
value CRYPT_STRING_NOCR (0x80000000)
value CRYPT_STRING_NOCRLF (0x40000000)
value CRYPT_STRING_PERCENTESCAPE (0x08000000)
value CRYPT_STRING_STRICT (0x20000000)
value CRYPT_SUCCEED (TRUE)
value CRYPT_TEMPLATE_OID_GROUP_ID (9)
value CRYPT_UI_PROMPT (0x00000004)
value CRYPT_UM ((0x00000001))
value CRYPT_UNICODE_NAME_ENCODE_DISABLE_CHECK_TYPE_FLAG (CERT_RDN_DISABLE_CHECK_TYPE_FLAG)
value CRYPT_UPDATE_KEY (0x00000008)
value CRYPT_USERDATA (1)
value CRYPT_USER_DEFAULT (0x00000002)
value CRYPT_USER_KEYSET (0x00001000)
value CRYPT_USER_PROTECTED (0x00000002)
value CRYPT_USER_PROTECTED_STRONG (0x00100000)
value CRYPT_VERIFYCONTEXT (0xF0000000)
value CRYPT_VERIFY_CERT_SIGN_CHECK_WEAK_HASH_FLAG (0x00000008)
value CRYPT_VERIFY_CERT_SIGN_ISSUER_CERT (2)
value CRYPT_VERIFY_CERT_SIGN_ISSUER_CHAIN (3)
value CRYPT_VERIFY_CERT_SIGN_ISSUER_NULL (4)
value CRYPT_VERIFY_CERT_SIGN_ISSUER_PUBKEY (1)
value CRYPT_VERIFY_CERT_SIGN_RETURN_STRONG_PROPERTIES_FLAG (0x00000004)
value CRYPT_VERIFY_CERT_SIGN_SET_STRONG_PROPERTIES_FLAG (0x00000002)
value CRYPT_VERIFY_CERT_SIGN_SUBJECT_BLOB (1)
value CRYPT_VERIFY_CERT_SIGN_SUBJECT_CERT (2)
value CRYPT_VERIFY_CERT_SIGN_SUBJECT_CRL (3)
value CRYPT_VERIFY_CERT_SIGN_SUBJECT_OCSP_BASIC_SIGNED_RESPONSE (4)
value CRYPT_VERIFY_CONTEXT_SIGNATURE (0x00000020)
value CRYPT_VERIFY_DATA_HASH (0x00000040)
value CRYPT_VOLATILE (0x00001000)
value CRYPT_WIRE_ONLY_RETRIEVAL (0x00000004)
value CRYPT_WRITE (0x0010)
value CRYPT_Y_ONLY (0x00000001)
value CSOUND_SYSTEM (16)
value CSTR_EQUAL (2)
value CSTR_GREATER_THAN (3)
value CSTR_LESS_THAN (1)
value CSV_INVALID_DEVICE_NUMBER (0xFFFFFFFF)
value CSV_MGMTLOCK_CHECK_VOLUME_REDIRECTED (0x00000001)
value CSV_QUERY_MDS_PATH_FLAG_CSV_DIRECT_IO_ENABLED (0x2)
value CSV_QUERY_MDS_PATH_FLAG_SMB_BYPASS_CSV_ENABLED (0x4)
value CSV_QUERY_MDS_PATH_FLAG_STORAGE_ON_THIS_NODE_IS_CONNECTED (0x1)
value CS_BYTEALIGNCLIENT (0x1000)
value CS_BYTEALIGNWINDOW (0x2000)
value CS_CLASSDC (0x0040)
value CS_DBLCLKS (0x0008)
value CS_DELETE_TRANSFORM (0x00000003L)
value CS_DISABLE (0x00000002L)
value CS_DROPSHADOW (0x00020000)
value CS_ENABLE (0x00000001L)
value CS_E_ADMIN_LIMIT_EXCEEDED (_HRESULT_TYPEDEF_(0x8004016DL))
value CS_E_CLASS_NOTFOUND (_HRESULT_TYPEDEF_(0x80040166L))
value CS_E_FIRST (0x80040164L)
value CS_E_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x8004016FL))
value CS_E_INVALID_PATH (_HRESULT_TYPEDEF_(0x8004016BL))
value CS_E_INVALID_VERSION (_HRESULT_TYPEDEF_(0x80040167L))
value CS_E_LAST (0x8004016FL)
value CS_E_NETWORK_ERROR (_HRESULT_TYPEDEF_(0x8004016CL))
value CS_E_NOT_DELETABLE (_HRESULT_TYPEDEF_(0x80040165L))
value CS_E_NO_CLASSSTORE (_HRESULT_TYPEDEF_(0x80040168L))
value CS_E_OBJECT_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x8004016AL))
value CS_E_OBJECT_NOTFOUND (_HRESULT_TYPEDEF_(0x80040169L))
value CS_E_PACKAGE_NOTFOUND (_HRESULT_TYPEDEF_(0x80040164L))
value CS_E_SCHEMA_MISMATCH (_HRESULT_TYPEDEF_(0x8004016EL))
value CS_GLOBALCLASS (0x4000)
value CS_HREDRAW (0x0002)
value CS_IME (0x00010000)
value CS_INSERTCHAR (0x2000)
value CS_NOCLOSE (0x0200)
value CS_NOMOVECARET (0x4000)
value CS_OWNDC (0x0020)
value CS_PARENTDC (0x0080)
value CS_SAVEBITS (0x0800)
value CS_VREDRAW (0x0001)
value CTLCOLOR_BTN (3)
value CTLCOLOR_DLG (4)
value CTLCOLOR_EDIT (1)
value CTLCOLOR_LISTBOX (2)
value CTLCOLOR_MAX (7)
value CTLCOLOR_MSGBOX (0)
value CTLCOLOR_SCROLLBAR (5)
value CTLCOLOR_STATIC (6)
value CTL_ANY_SUBJECT_TYPE (1)
value CTL_CERT_SUBJECT_TYPE (2)
value CTL_ENTRY_FROM_PROP_CHAIN_FLAG (0x1)
value CTL_FIND_ANY (0)
value CTL_FIND_EXISTING (5)
value CTL_FIND_NO_LIST_ID_CBDATA (0xFFFFFFFF)
value CTL_FIND_NO_SIGNER_PTR (((PCERT_INFO) -1))
value CTL_FIND_SAME_USAGE_FLAG (0x1)
value CTL_FIND_SUBJECT (4)
value CTL_FIND_USAGE (3)
value CTMF_INCLUDE_APPCONTAINER (0x00000001UL)
value CTMF_INCLUDE_LPAC (0x00000002UL)
value CTMF_VALID_FLAGS ((CTMF_INCLUDE_APPCONTAINER | CTMF_INCLUDE_LPAC))
value CTRL_BREAK_EVENT (1)
value CTRL_CLOSE_EVENT (2)
value CTRL_C_EVENT (0)
value CTRL_LOGOFF_EVENT (5)
value CTRL_SHUTDOWN_EVENT (6)
value CTRY_ALBANIA (355)
value CTRY_ALGERIA (213)
value CTRY_ARGENTINA (54)
value CTRY_ARMENIA (374)
value CTRY_AUSTRALIA (61)
value CTRY_AUSTRIA (43)
value CTRY_AZERBAIJAN (994)
value CTRY_BAHRAIN (973)
value CTRY_BELARUS (375)
value CTRY_BELGIUM (32)
value CTRY_BELIZE (501)
value CTRY_BOLIVIA (591)
value CTRY_BRAZIL (55)
value CTRY_BRUNEI_DARUSSALAM (673)
value CTRY_BULGARIA (359)
value CTRY_CANADA (2)
value CTRY_CARIBBEAN (1)
value CTRY_CHILE (56)
value CTRY_COLOMBIA (57)
value CTRY_COSTA_RICA (506)
value CTRY_CROATIA (385)
value CTRY_CZECH (420)
value CTRY_DEFAULT (0)
value CTRY_DENMARK (45)
value CTRY_DOMINICAN_REPUBLIC (1)
value CTRY_ECUADOR (593)
value CTRY_EGYPT (20)
value CTRY_EL_SALVADOR (503)
value CTRY_ESTONIA (372)
value CTRY_FAEROE_ISLANDS (298)
value CTRY_FINLAND (358)
value CTRY_FRANCE (33)
value CTRY_GEORGIA (995)
value CTRY_GERMANY (49)
value CTRY_GREECE (30)
value CTRY_GUATEMALA (502)
value CTRY_HONDURAS (504)
value CTRY_HONG_KONG (852)
value CTRY_HUNGARY (36)
value CTRY_ICELAND (354)
value CTRY_INDIA (91)
value CTRY_INDONESIA (62)
value CTRY_IRAN (981)
value CTRY_IRAQ (964)
value CTRY_IRELAND (353)
value CTRY_ISRAEL (972)
value CTRY_ITALY (39)
value CTRY_JAMAICA (1)
value CTRY_JAPAN (81)
value CTRY_JORDAN (962)
value CTRY_KAZAKSTAN (7)
value CTRY_KENYA (254)
value CTRY_KUWAIT (965)
value CTRY_KYRGYZSTAN (996)
value CTRY_LATVIA (371)
value CTRY_LEBANON (961)
value CTRY_LIBYA (218)
value CTRY_LIECHTENSTEIN (41)
value CTRY_LITHUANIA (370)
value CTRY_LUXEMBOURG (352)
value CTRY_MACAU (853)
value CTRY_MACEDONIA (389)
value CTRY_MALAYSIA (60)
value CTRY_MALDIVES (960)
value CTRY_MEXICO (52)
value CTRY_MONACO (33)
value CTRY_MONGOLIA (976)
value CTRY_MOROCCO (212)
value CTRY_NETHERLANDS (31)
value CTRY_NEW_ZEALAND (64)
value CTRY_NICARAGUA (505)
value CTRY_NORWAY (47)
value CTRY_OMAN (968)
value CTRY_PAKISTAN (92)
value CTRY_PANAMA (507)
value CTRY_PARAGUAY (595)
value CTRY_PERU (51)
value CTRY_PHILIPPINES (63)
value CTRY_POLAND (48)
value CTRY_PORTUGAL (351)
value CTRY_PRCHINA (86)
value CTRY_PUERTO_RICO (1)
value CTRY_QATAR (974)
value CTRY_ROMANIA (40)
value CTRY_RUSSIA (7)
value CTRY_SAUDI_ARABIA (966)
value CTRY_SERBIA (381)
value CTRY_SINGAPORE (65)
value CTRY_SLOVAK (421)
value CTRY_SLOVENIA (386)
value CTRY_SOUTH_AFRICA (27)
value CTRY_SOUTH_KOREA (82)
value CTRY_SPAIN (34)
value CTRY_SWEDEN (46)
value CTRY_SWITZERLAND (41)
value CTRY_SYRIA (963)
value CTRY_TAIWAN (886)
value CTRY_TATARSTAN (7)
value CTRY_THAILAND (66)
value CTRY_TRINIDAD_Y_TOBAGO (1)
value CTRY_TUNISIA (216)
value CTRY_TURKEY (90)
value CTRY_UAE (971)
value CTRY_UKRAINE (380)
value CTRY_UNITED_KINGDOM (44)
value CTRY_UNITED_STATES (1)
value CTRY_URUGUAY (598)
value CTRY_UZBEKISTAN (7)
value CTRY_VENEZUELA (58)
value CTRY_VIET_NAM (84)
value CTRY_YEMEN (967)
value CTRY_ZIMBABWE (263)
value CURRENT_IMPORT_REDIRECTION_VERSION (1)
value CURSOR_CREATION_SCALING_DEFAULT (2)
value CURSOR_CREATION_SCALING_NONE (1)
value CURSOR_SHOWING (0x00000001)
value CURSOR_SUPPRESSED (0x00000002)
value CURVECAPS (28)
value CUR_BLOB_VERSION (2)
value CWCSTORAGENAME (32)
value CWF_CREATE_ONLY (0x00000001)
value CWMO_MAX_HANDLES (56)
value CWP_ALL (0x0000)
value CWP_SKIPDISABLED (0x0002)
value CWP_SKIPINVISIBLE (0x0001)
value CWP_SKIPTRANSPARENT (0x0004)
value DACL_SECURITY_INFORMATION ((0x00000004L))
value DATA_E_FIRST (0x80040130L)
value DATA_E_FORMATETC (DV_E_FORMATETC)
value DATA_E_LAST (0x8004013FL)
value DATA_S_FIRST (0x00040130L)
value DATA_S_LAST (0x0004013FL)
value DATA_S_SAMEFORMATETC (_HRESULT_TYPEDEF_(0x00040130L))
value DATEFMT_ENUMPROC (DATEFMT_ENUMPROCA)
value DATEFMT_ENUMPROCEX (DATEFMT_ENUMPROCEXA)
value DATE_AUTOLAYOUT (0x00000040)
value DATE_LONGDATE (0x00000002)
value DATE_LTRREADING (0x00000010)
value DATE_MONTHDAY (0x00000080)
value DATE_RTLREADING (0x00000020)
value DATE_SHORTDATE (0x00000001)
value DATE_USE_ALT_CALENDAR (0x00000004)
value DATE_YEARMONTH (0x00000008)
value DAX_ALLOC_ALIGNMENT_FLAG_FALLBACK_SPECIFIED ((0x00000002))
value DAX_ALLOC_ALIGNMENT_FLAG_MANDATORY ((0x00000001))
value DBG_COMMAND_EXCEPTION (((DWORD )0x40010009L))
value DBG_CONTINUE (((DWORD )0x00010002L))
value DBG_CONTROL_BREAK (((DWORD )0x40010008L))
value DBG_CONTROL_C (((DWORD )0x40010005L))
value DBG_EXCEPTION_HANDLED (((DWORD )0x00010001L))
value DBG_EXCEPTION_NOT_HANDLED (((DWORD )0x80010001L))
value DBG_PRINTEXCEPTION_C (((DWORD )0x40010006L))
value DBG_PRINTEXCEPTION_WIDE_C (((DWORD )0x4001000AL))
value DBG_REPLY_LATER (((DWORD )0x40010001L))
value DBG_RIPEXCEPTION (((DWORD )0x40010007L))
value DBG_TERMINATE_PROCESS (((DWORD )0x40010004L))
value DBG_TERMINATE_THREAD (((DWORD )0x40010003L))
value DCBA_FACEDOWNCENTER (0x0101)
value DCBA_FACEDOWNLEFT (0x0102)
value DCBA_FACEDOWNNONE (0x0100)
value DCBA_FACEDOWNRIGHT (0x0103)
value DCBA_FACEUPCENTER (0x0001)
value DCBA_FACEUPLEFT (0x0002)
value DCBA_FACEUPNONE (0x0000)
value DCBA_FACEUPRIGHT (0x0003)
value DCB_ACCUMULATE (0x0002)
value DCB_DIRTY (DCB_ACCUMULATE)
value DCB_DISABLE (0x0008)
value DCB_ENABLE (0x0004)
value DCB_RESET (0x0001)
value DCB_SET ((DCB_RESET | DCB_ACCUMULATE))
value DCE_C_ERROR_STRING_LEN (256)
value DCOMPOSITION_ERROR_SURFACE_BEING_RENDERED (_HRESULT_TYPEDEF_(0x88980801L))
value DCOMPOSITION_ERROR_SURFACE_NOT_BEING_RENDERED (_HRESULT_TYPEDEF_(0x88980802L))
value DCOMPOSITION_ERROR_WINDOW_ALREADY_COMPOSED (_HRESULT_TYPEDEF_(0x88980800L))
value DCOMSCM_ACTIVATION_DISALLOW_UNSECURE_CALL (0x2)
value DCOMSCM_ACTIVATION_USE_ALL_AUTHNSERVICES (0x1)
value DCOMSCM_PING_DISALLOW_UNSECURE_CALL (0x20)
value DCOMSCM_PING_USE_MID_AUTHNSERVICE (0x10)
value DCOMSCM_RESOLVE_DISALLOW_UNSECURE_CALL (0x8)
value DCOMSCM_RESOLVE_USE_ALL_AUTHNSERVICES (0x4)
value DCTT_BITMAP (0x0000001L)
value DCTT_DOWNLOAD (0x0000002L)
value DCTT_DOWNLOAD_OUTLINE (0x0000008L)
value DCTT_SUBDEV (0x0000004L)
value DCX_CACHE (0x00000002L)
value DCX_CLIPCHILDREN (0x00000008L)
value DCX_CLIPSIBLINGS (0x00000010L)
value DCX_EXCLUDERGN (0x00000040L)
value DCX_EXCLUDEUPDATE (0x00000100L)
value DCX_INTERSECTRGN (0x00000080L)
value DCX_INTERSECTUPDATE (0x00000200L)
value DCX_LOCKWINDOWUPDATE (0x00000400L)
value DCX_NORESETATTRS (0x00000004L)
value DCX_PARENTCLIP (0x00000020L)
value DCX_VALIDATE (0x00200000L)
value DCX_WINDOW (0x00000001L)
value DC_ACTIVE (0x0001)
value DC_BINADJUST (19)
value DC_BINNAMES (12)
value DC_BINS (6)
value DC_BRUSH (18)
value DC_BUTTONS (0x1000)
value DC_COLLATE (22)
value DC_COLORDEVICE (32)
value DC_COPIES (18)
value DC_DATATYPE_PRODUCED (21)
value DC_DRIVER (11)
value DC_DUPLEX (7)
value DC_EMF_COMPLIANT (20)
value DC_ENUMRESOLUTIONS (13)
value DC_EXTRA (9)
value DC_FIELDS (1)
value DC_FILEDEPENDENCIES (14)
value DC_GRADIENT (0x0020)
value DC_HASDEFID (0x534B)
value DC_ICON (0x0004)
value DC_INBUTTON (0x0010)
value DC_MANUFACTURER (23)
value DC_MAXEXTENT (5)
value DC_MEDIAREADY (29)
value DC_MEDIATYPENAMES (34)
value DC_MEDIATYPES (35)
value DC_MINEXTENT (4)
value DC_MODEL (24)
value DC_NUP (33)
value DC_ORIENTATION (17)
value DC_PAPERNAMES (16)
value DC_PAPERS (2)
value DC_PAPERSIZE (3)
value DC_PEN (19)
value DC_PERSONALITY (25)
value DC_PRINTERMEM (28)
value DC_PRINTRATE (26)
value DC_PRINTRATEPPM (31)
value DC_PRINTRATEUNIT (27)
value DC_SIZE (8)
value DC_SMALLCAP (0x0002)
value DC_STAPLE (30)
value DC_TEXT (0x0008)
value DC_TRUETYPE (15)
value DC_VERSION (10)
value DDD_EXACT_MATCH_ON_REMOVE (0x00000004)
value DDD_LUID_BROADCAST_DRIVE (0x00000010)
value DDD_NO_BROADCAST_SYSTEM (0x00000008)
value DDD_RAW_TARGET_PATH (0x00000001)
value DDD_REMOVE_DEFINITION (0x00000002)
value DDE_FACK (0x8000)
value DDE_FACKREQ (0x8000)
value DDE_FAPPSTATUS (0x00ff)
value DDE_FBUSY (0x4000)
value DDE_FDEFERUPD (0x4000)
value DDE_FNOTPROCESSED (0x0000)
value DDE_FRELEASE (0x2000)
value DDE_FREQUESTED (0x1000)
value DDL_ARCHIVE (0x0020)
value DDL_DIRECTORY (0x0010)
value DDL_DRIVES (0x4000)
value DDL_EXCLUSIVE (0x8000)
value DDL_HIDDEN (0x0002)
value DDL_POSTMSGS (0x2000)
value DDL_READONLY (0x0001)
value DDL_READWRITE (0x0000)
value DDL_SYSTEM (0x0004)
value DDUMP_FLAG_DATA_READ_FROM_DEVICE (0x0001)
value DD_DEFDRAGDELAY (( 200 ))
value DD_DEFDRAGMINDIST (( 2 ))
value DD_DEFSCROLLDELAY (( 50 ))
value DD_DEFSCROLLINSET (( 11 ))
value DD_DEFSCROLLINTERVAL (( 50 ))
value DEACTIVATE_ACTCTX_FLAG_FORCE_EARLY_DEACTIVATION ((0x00000001))
value DEBUG_ONLY_THIS_PROCESS (0x00000002)
value DEBUG_PROCESS (0x00000001)
value DECIMAL_NEG (((BYTE)0x80))
value DECLSPEC_CACHEALIGN (DECLSPEC_ALIGN(SYSTEM_CACHE_ALIGNMENT_SIZE))
value DEDICATED_MEMORY_CACHE_ELIGIBLE (0x1)
value DEFAULT_CHARSET (1)
value DEFAULT_GUI_FONT (17)
value DEFAULT_PALETTE (15)
value DEFAULT_PITCH (0)
value DEFAULT_QUALITY (0)
value DEF_PRIORITY (1)
value DELETE ((0x00010000L))
value DEREGISTERED (0x05)
value DESKTOPHORZRES (118)
value DESKTOPVERTRES (117)
value DESKTOP_CREATEMENU (0x0004L)
value DESKTOP_CREATEWINDOW (0x0002L)
value DESKTOP_ENUMERATE (0x0040L)
value DESKTOP_HOOKCONTROL (0x0008L)
value DESKTOP_JOURNALPLAYBACK (0x0020L)
value DESKTOP_JOURNALRECORD (0x0010L)
value DESKTOP_READOBJECTS (0x0001L)
value DESKTOP_SWITCHDESKTOP (0x0100L)
value DESKTOP_WRITEOBJECTS (0x0080L)
value DETACHED_PROCESS (0x00000008)
value DEVICEDATA (19)
value DEVICEDUMP_CAP_PRIVATE_SECTION (0x00000001)
value DEVICEDUMP_CAP_RESTRICTED_SECTION (0x00000002)
value DEVICEDUMP_MAX_IDSTRING (32)
value DEVICEFAMILYDEVICEFORM_ALLINONE (0x00000007)
value DEVICEFAMILYDEVICEFORM_BANKING (0x0000000E)
value DEVICEFAMILYDEVICEFORM_BUILDING_AUTOMATION (0x0000000F)
value DEVICEFAMILYDEVICEFORM_CONVERTIBLE (0x00000005)
value DEVICEFAMILYDEVICEFORM_DESKTOP (0x00000003)
value DEVICEFAMILYDEVICEFORM_DETACHABLE (0x00000006)
value DEVICEFAMILYDEVICEFORM_DIGITAL_SIGNAGE (0x00000010)
value DEVICEFAMILYDEVICEFORM_GAMING (0x00000011)
value DEVICEFAMILYDEVICEFORM_HMD (0x0000000B)
value DEVICEFAMILYDEVICEFORM_HOME_AUTOMATION (0x00000012)
value DEVICEFAMILYDEVICEFORM_INDUSTRIAL_AUTOMATION (0x00000013)
value DEVICEFAMILYDEVICEFORM_INDUSTRY_HANDHELD (0x0000000C)
value DEVICEFAMILYDEVICEFORM_INDUSTRY_OTHER (0x0000001D)
value DEVICEFAMILYDEVICEFORM_INDUSTRY_TABLET (0x0000000D)
value DEVICEFAMILYDEVICEFORM_KIOSK (0x00000014)
value DEVICEFAMILYDEVICEFORM_LARGESCREEN (0x0000000A)
value DEVICEFAMILYDEVICEFORM_MAKER_BOARD (0x00000015)
value DEVICEFAMILYDEVICEFORM_MAX (0x0000002D)
value DEVICEFAMILYDEVICEFORM_MEDICAL (0x00000016)
value DEVICEFAMILYDEVICEFORM_NETWORKING (0x00000017)
value DEVICEFAMILYDEVICEFORM_NOTEBOOK (0x00000004)
value DEVICEFAMILYDEVICEFORM_PHONE (0x00000001)
value DEVICEFAMILYDEVICEFORM_POINT_OF_SERVICE (0x00000018)
value DEVICEFAMILYDEVICEFORM_PRINTING (0x00000019)
value DEVICEFAMILYDEVICEFORM_PUCK (0x00000009)
value DEVICEFAMILYDEVICEFORM_STICKPC (0x00000008)
value DEVICEFAMILYDEVICEFORM_TABLET (0x00000002)
value DEVICEFAMILYDEVICEFORM_THIN_CLIENT (0x0000001A)
value DEVICEFAMILYDEVICEFORM_TOY (0x0000001B)
value DEVICEFAMILYDEVICEFORM_UNKNOWN (0x00000000)
value DEVICEFAMILYDEVICEFORM_VENDING (0x0000001C)
value DEVICEFAMILYDEVICEFORM_XBOX_ONE (0x0000001E)
value DEVICEFAMILYDEVICEFORM_XBOX_ONE_S (0x0000001F)
value DEVICEFAMILYDEVICEFORM_XBOX_ONE_X (0x00000020)
value DEVICEFAMILYDEVICEFORM_XBOX_ONE_X_DEVKIT (0x00000021)
value DEVICEFAMILYDEVICEFORM_XBOX_SERIES_S (0x00000024)
value DEVICEFAMILYDEVICEFORM_XBOX_SERIES_X (0x00000022)
value DEVICEFAMILYDEVICEFORM_XBOX_SERIES_X_DEVKIT (0x00000023)
value DEVICEFAMILYINFOENUM_DESKTOP (0x00000003)
value DEVICEFAMILYINFOENUM_HOLOGRAPHIC (0x0000000A)
value DEVICEFAMILYINFOENUM_IOT (0x00000007)
value DEVICEFAMILYINFOENUM_IOT_HEADLESS (0x00000008)
value DEVICEFAMILYINFOENUM_MAX (0x00000011)
value DEVICEFAMILYINFOENUM_MOBILE (0x00000004)
value DEVICEFAMILYINFOENUM_SERVER (0x00000009)
value DEVICEFAMILYINFOENUM_SERVER_NANO (0x0000000D)
value DEVICEFAMILYINFOENUM_TEAM (0x00000006)
value DEVICEFAMILYINFOENUM_UAP (0x00000000)
value DEVICEFAMILYINFOENUM_WINDOWS_CORE (0x00000010)
value DEVICEFAMILYINFOENUM_WINDOWS_CORE_HEADLESS (0x00000011)
value DEVICEFAMILYINFOENUM_XBOX (0x00000005)
value DEVICEFAMILYINFOENUM_XBOXERA (0x0000000C)
value DEVICEFAMILYINFOENUM_XBOXSRA (0x0000000B)
value DEVICE_DEFAULT_FONT (14)
value DEVICE_DSM_FLAG_ALLOCATION_CONSOLIDATEABLE_ONLY (0x40000000)
value DEVICE_DSM_FLAG_ENTIRE_DATA_SET_RANGE (0x00000001)
value DEVICE_DSM_FLAG_PHYSICAL_ADDRESSES_OMIT_TOTAL_RANGES (0x10000000)
value DEVICE_DSM_FLAG_REPAIR_INPUT_TOPOLOGY_ID_PRESENT (0x40000000)
value DEVICE_DSM_FLAG_REPAIR_OUTPUT_PARITY_EXTENT (0x20000000)
value DEVICE_DSM_FLAG_SCRUB_OUTPUT_PARITY_EXTENT (0x20000000)
value DEVICE_DSM_FLAG_SCRUB_SKIP_IN_SYNC (0x10000000)
value DEVICE_DSM_FLAG_TRIM_BYPASS_RZAT (0x40000000)
value DEVICE_DSM_FLAG_TRIM_NOT_FS_ALLOCATED (0x80000000)
value DEVICE_DSM_NOTIFY_FLAG_BEGIN (0x00000001)
value DEVICE_DSM_NOTIFY_FLAG_END (0x00000002)
value DEVICE_DSM_PHYSICAL_ADDRESS_HAS_MEMORY_ERROR (((LONGLONG)-1))
value DEVICE_FONTTYPE (0x0002)
value DEVICE_NOTIFY_ALL_INTERFACE_CLASSES (0x00000004)
value DEVICE_NOTIFY_SERVICE_HANDLE (0x00000001)
value DEVICE_NOTIFY_WINDOW_HANDLE (0x00000000)
value DEVICE_STORAGE_NO_ERRORS (0x1)
value DEVICE_TYPE (DWORD)
value DFCS_ADJUSTRECT (0x2000)
value DFCS_BUTTONCHECK (0x0000)
value DFCS_BUTTONPUSH (0x0010)
value DFCS_BUTTONRADIO (0x0004)
value DFCS_BUTTONRADIOIMAGE (0x0001)
value DFCS_BUTTONRADIOMASK (0x0002)
value DFCS_CAPTIONCLOSE (0x0000)
value DFCS_CAPTIONHELP (0x0004)
value DFCS_CAPTIONMAX (0x0002)
value DFCS_CAPTIONMIN (0x0001)
value DFCS_CAPTIONRESTORE (0x0003)
value DFCS_CHECKED (0x0400)
value DFCS_FLAT (0x4000)
value DFCS_HOT (0x1000)
value DFCS_INACTIVE (0x0100)
value DFCS_MENUARROW (0x0000)
value DFCS_MENUARROWRIGHT (0x0004)
value DFCS_MENUBULLET (0x0002)
value DFCS_MENUCHECK (0x0001)
value DFCS_MONO (0x8000)
value DFCS_PUSHED (0x0200)
value DFCS_SCROLLCOMBOBOX (0x0005)
value DFCS_SCROLLDOWN (0x0001)
value DFCS_SCROLLLEFT (0x0002)
value DFCS_SCROLLRIGHT (0x0003)
value DFCS_SCROLLSIZEGRIP (0x0008)
value DFCS_SCROLLSIZEGRIPRIGHT (0x0010)
value DFCS_SCROLLUP (0x0000)
value DFCS_TRANSPARENT (0x0800)
value DFC_BUTTON (4)
value DFC_CAPTION (1)
value DFC_MENU (2)
value DFC_POPUPMENU (5)
value DFC_SCROLL (3)
value DF_ALLOWOTHERACCOUNTHOOK (0x0001L)
value DIAGNOSTIC_REASON_DETAILED_STRING (0x00000002)
value DIAGNOSTIC_REASON_NOT_SPECIFIED (0x80000000)
value DIAGNOSTIC_REASON_SIMPLE_STRING (0x00000001)
value DIAGNOSTIC_REASON_VERSION (0)
value DIALOPTION_BILLING (0x00000040)
value DIALOPTION_DIALTONE (0x00000100)
value DIALOPTION_QUIET (0x00000080)
value DIB_PAL_COLORS (1)
value DIB_RGB_COLORS (0)
value DIFFERENCE (11)
value DIGSIG_E_CRYPTO (_HRESULT_TYPEDEF_(0x800B0008L))
value DIGSIG_E_DECODE (_HRESULT_TYPEDEF_(0x800B0006L))
value DIGSIG_E_ENCODE (_HRESULT_TYPEDEF_(0x800B0005L))
value DIGSIG_E_EXTENSIBILITY (_HRESULT_TYPEDEF_(0x800B0007L))
value DISABLE_MAX_PRIVILEGE (0x1)
value DISABLE_NEWLINE_AUTO_RETURN (0x0008)
value DISABLE_SMART (0xD9)
value DISCHARGE_POLICY_CRITICAL (0)
value DISCHARGE_POLICY_LOW (1)
value DISC_NO_FORCE (0x00000040)
value DISC_UPDATE_PROFILE (0x00000001)
value DISK_ATTRIBUTE_OFFLINE (0x0000000000000001)
value DISK_ATTRIBUTE_READ_ONLY (0x0000000000000002)
value DISK_BINNING (3)
value DISK_LOGGING_DUMP (2)
value DISK_LOGGING_START (0)
value DISK_LOGGING_STOP (1)
value DISPATCH_LEVEL (2)
value DISPATCH_METHOD (0x1)
value DISPATCH_PROPERTYGET (0x2)
value DISPATCH_PROPERTYPUT (0x4)
value DISPATCH_PROPERTYPUTREF (0x8)
value DISPID_COLLECT (( -8 ))
value DISPID_CONSTRUCTOR (( -6 ))
value DISPID_DESTRUCTOR (( -7 ))
value DISPID_EVALUATE (( -5 ))
value DISPID_NEWENUM (( -4 ))
value DISPID_PROPERTYPUT (( -3 ))
value DISPID_UNKNOWN (( -1 ))
value DISPID_VALUE (( 0 ))
value DISPLAYCONFIG_MAXPATH (1024)
value DISPLAYCONFIG_PATH_ACTIVE (0x00000001)
value DISPLAYCONFIG_PATH_CLONE_GROUP_INVALID (0xffff)
value DISPLAYCONFIG_PATH_DESKTOP_IMAGE_IDX_INVALID (0xffff)
value DISPLAYCONFIG_PATH_MODE_IDX_INVALID (0xffffffff)
value DISPLAYCONFIG_PATH_PREFERRED_UNSCALED (0x00000004)
value DISPLAYCONFIG_PATH_SOURCE_MODE_IDX_INVALID (0xffff)
value DISPLAYCONFIG_PATH_SUPPORT_VIRTUAL_MODE (0x00000008)
value DISPLAYCONFIG_PATH_TARGET_MODE_IDX_INVALID (0xffff)
value DISPLAYCONFIG_PATH_VALID_FLAGS (0x0000001D)
value DISPLAYCONFIG_SOURCE_IN_USE (0x00000001)
value DISPLAYCONFIG_TARGET_FORCED_AVAILABILITY_BOOT (0x00000004)
value DISPLAYCONFIG_TARGET_FORCED_AVAILABILITY_PATH (0x00000008)
value DISPLAYCONFIG_TARGET_FORCED_AVAILABILITY_SYSTEM (0x00000010)
value DISPLAYCONFIG_TARGET_FORCIBLE (0x00000002)
value DISPLAYCONFIG_TARGET_IN_USE (0x00000001)
value DISPLAYCONFIG_TARGET_IS_HMD (0x00000020)
value DISPLAY_DEVICE_ACC_DRIVER (0x00000040)
value DISPLAY_DEVICE_ACTIVE (0x00000001)
value DISPLAY_DEVICE_ATTACHED (0x00000002)
value DISPLAY_DEVICE_ATTACHED_TO_DESKTOP (0x00000001)
value DISPLAY_DEVICE_DISCONNECT (0x02000000)
value DISPLAY_DEVICE_MIRRORING_DRIVER (0x00000008)
value DISPLAY_DEVICE_MODESPRUNED (0x08000000)
value DISPLAY_DEVICE_MULTI_DRIVER (0x00000002)
value DISPLAY_DEVICE_PRIMARY_DEVICE (0x00000004)
value DISPLAY_DEVICE_RDPUDD (0x01000000)
value DISPLAY_DEVICE_REMOTE (0x04000000)
value DISPLAY_DEVICE_REMOVABLE (0x00000020)
value DISPLAY_DEVICE_TS_COMPATIBLE (0x00200000)
value DISPLAY_DEVICE_UNSAFE_MODES_ON (0x00080000)
value DISPLAY_DEVICE_VGA_COMPATIBLE (0x00000010)
value DISP_CHANGE_BADDUALVIEW (-6)
value DISP_CHANGE_BADFLAGS (-4)
value DISP_CHANGE_BADMODE (-2)
value DISP_CHANGE_BADPARAM (-5)
value DISP_CHANGE_FAILED (-1)
value DISP_CHANGE_NOTUPDATED (-3)
value DISP_CHANGE_RESTART (1)
value DISP_CHANGE_SUCCESSFUL (0)
value DISP_E_ARRAYISLOCKED (_HRESULT_TYPEDEF_(0x8002000DL))
value DISP_E_BADCALLEE (_HRESULT_TYPEDEF_(0x80020010L))
value DISP_E_BADINDEX (_HRESULT_TYPEDEF_(0x8002000BL))
value DISP_E_BADPARAMCOUNT (_HRESULT_TYPEDEF_(0x8002000EL))
value DISP_E_BADVARTYPE (_HRESULT_TYPEDEF_(0x80020008L))
value DISP_E_BUFFERTOOSMALL (_HRESULT_TYPEDEF_(0x80020013L))
value DISP_E_DIVBYZERO (_HRESULT_TYPEDEF_(0x80020012L))
value DISP_E_EXCEPTION (_HRESULT_TYPEDEF_(0x80020009L))
value DISP_E_MEMBERNOTFOUND (_HRESULT_TYPEDEF_(0x80020003L))
value DISP_E_NONAMEDARGS (_HRESULT_TYPEDEF_(0x80020007L))
value DISP_E_NOTACOLLECTION (_HRESULT_TYPEDEF_(0x80020011L))
value DISP_E_OVERFLOW (_HRESULT_TYPEDEF_(0x8002000AL))
value DISP_E_PARAMNOTFOUND (_HRESULT_TYPEDEF_(0x80020004L))
value DISP_E_PARAMNOTOPTIONAL (_HRESULT_TYPEDEF_(0x8002000FL))
value DISP_E_TYPEMISMATCH (_HRESULT_TYPEDEF_(0x80020005L))
value DISP_E_UNKNOWNINTERFACE (_HRESULT_TYPEDEF_(0x80020001L))
value DISP_E_UNKNOWNLCID (_HRESULT_TYPEDEF_(0x8002000CL))
value DISP_E_UNKNOWNNAME (_HRESULT_TYPEDEF_(0x80020006L))
value DI_APPBANDING (0x00000001)
value DI_CHANNEL (1)
value DI_COMPAT (0x0004)
value DI_DEFAULTSIZE (0x0008)
value DI_IMAGE (0x0002)
value DI_MASK (0x0001)
value DI_MEMORYMAP_WRITE (0x00000001)
value DI_NOMIRROR (0x0010)
value DI_NORMAL (0x0003)
value DI_READ_SPOOL_JOB (3)
value DI_ROPS_READ_DESTINATION (0x00000002)
value DKGRAY_BRUSH (3)
value DLGC_BUTTON (0x2000)
value DLGC_DEFPUSHBUTTON (0x0010)
value DLGC_HASSETSEL (0x0008)
value DLGC_RADIOBUTTON (0x0040)
value DLGC_STATIC (0x0100)
value DLGC_UNDEFPUSHBUTTON (0x0020)
value DLGC_WANTALLKEYS (0x0004)
value DLGC_WANTARROWS (0x0001)
value DLGC_WANTCHARS (0x0080)
value DLGC_WANTMESSAGE (0x0004)
value DLGC_WANTTAB (0x0002)
value DLGWINDOWEXTRA (30)
value DLL_PROCESS_ATTACH (1)
value DLL_PROCESS_DETACH (0)
value DLL_THREAD_ATTACH (2)
value DLL_THREAD_DETACH (3)
value DMBIN_AUTO (7)
value DMBIN_CASSETTE (14)
value DMBIN_ENVELOPE (5)
value DMBIN_ENVMANUAL (6)
value DMBIN_FIRST (DMBIN_UPPER)
value DMBIN_FORMSOURCE (15)
value DMBIN_LARGECAPACITY (11)
value DMBIN_LARGEFMT (10)
value DMBIN_LAST (DMBIN_FORMSOURCE)
value DMBIN_LOWER (2)
value DMBIN_MANUAL (4)
value DMBIN_MIDDLE (3)
value DMBIN_ONLYONE (1)
value DMBIN_SMALLFMT (9)
value DMBIN_TRACTOR (8)
value DMBIN_UPPER (1)
value DMBIN_USER (256)
value DMCOLLATE_FALSE (0)
value DMCOLLATE_TRUE (1)
value DMCOLOR_COLOR (2)
value DMCOLOR_MONOCHROME (1)
value DMDFO_CENTER (2)
value DMDFO_DEFAULT (0)
value DMDFO_STRETCH (1)
value DMDISPLAYFLAGS_TEXTMODE (0x00000004)
value DMDITHER_COARSE (2)
value DMDITHER_ERRORDIFFUSION (5)
value DMDITHER_FINE (3)
value DMDITHER_GRAYSCALE (10)
value DMDITHER_LINEART (4)
value DMDITHER_NONE (1)
value DMDITHER_USER (256)
value DMDO_DEFAULT (0)
value DMDUP_HORIZONTAL (3)
value DMDUP_SIMPLEX (1)
value DMDUP_VERTICAL (2)
value DMICMMETHOD_DEVICE (4)
value DMICMMETHOD_DRIVER (3)
value DMICMMETHOD_NONE (1)
value DMICMMETHOD_SYSTEM (2)
value DMICMMETHOD_USER (256)
value DMICM_ABS_COLORIMETRIC (4)
value DMICM_COLORIMETRIC (3)
value DMICM_CONTRAST (2)
value DMICM_SATURATE (1)
value DMICM_USER (256)
value DMLERR_ADVACKTIMEOUT (0x4000)
value DMLERR_BUSY (0x4001)
value DMLERR_DATAACKTIMEOUT (0x4002)
value DMLERR_DLL_NOT_INITIALIZED (0x4003)
value DMLERR_DLL_USAGE (0x4004)
value DMLERR_EXECACKTIMEOUT (0x4005)
value DMLERR_FIRST (0x4000)
value DMLERR_INVALIDPARAMETER (0x4006)
value DMLERR_LAST (0x4011)
value DMLERR_LOW_MEMORY (0x4007)
value DMLERR_MEMORY_ERROR (0x4008)
value DMLERR_NOTPROCESSED (0x4009)
value DMLERR_NO_CONV_ESTABLISHED (0x400a)
value DMLERR_NO_ERROR (0)
value DMLERR_POKEACKTIMEOUT (0x400b)
value DMLERR_POSTMSG_FAILED (0x400c)
value DMLERR_REENTRANCY (0x400d)
value DMLERR_SERVER_DIED (0x400e)
value DMLERR_SYS_ERROR (0x400f)
value DMLERR_UNADVACKTIMEOUT (0x4010)
value DMLERR_UNFOUND_QUEUE_ID (0x4011)
value DMMEDIA_GLOSSY (3)
value DMMEDIA_STANDARD (1)
value DMMEDIA_TRANSPARENCY (2)
value DMMEDIA_USER (256)
value DMNUP_ONEUP (2)
value DMNUP_SYSTEM (1)
value DMORIENT_LANDSCAPE (2)
value DMORIENT_PORTRAIT (1)
value DMPAPER_A_PLUS (57)
value DMPAPER_B_PLUS (58)
value DMPAPER_CSHEET (24)
value DMPAPER_DBL_JAPANESE_POSTCARD (69)
value DMPAPER_DBL_JAPANESE_POSTCARD_ROTATED (82)
value DMPAPER_DSHEET (25)
value DMPAPER_ENV_DL (27)
value DMPAPER_ENV_INVITE (47)
value DMPAPER_ENV_ITALY (36)
value DMPAPER_ENV_MONARCH (37)
value DMPAPER_ENV_PERSONAL (38)
value DMPAPER_ESHEET (26)
value DMPAPER_EXECUTIVE (7)
value DMPAPER_FANFOLD_LGL_GERMAN (41)
value DMPAPER_FANFOLD_STD_GERMAN (40)
value DMPAPER_FANFOLD_US (39)
value DMPAPER_FIRST (DMPAPER_LETTER)
value DMPAPER_FOLIO (14)
value DMPAPER_JAPANESE_POSTCARD (43)
value DMPAPER_JAPANESE_POSTCARD_ROTATED (81)
value DMPAPER_LAST (DMPAPER_PENV_10_ROTATED)
value DMPAPER_LEDGER (4)
value DMPAPER_LEGAL (5)
value DMPAPER_LEGAL_EXTRA (51)
value DMPAPER_LETTER (1)
value DMPAPER_LETTERSMALL (2)
value DMPAPER_LETTER_EXTRA (50)
value DMPAPER_LETTER_EXTRA_TRANSVERSE (56)
value DMPAPER_LETTER_PLUS (59)
value DMPAPER_LETTER_ROTATED (75)
value DMPAPER_LETTER_TRANSVERSE (54)
value DMPAPER_NOTE (18)
value DMPAPER_QUARTO (15)
value DMPAPER_STATEMENT (6)
value DMPAPER_TABLOID (3)
value DMPAPER_TABLOID_EXTRA (52)
value DMPAPER_USER (256)
value DMRES_DRAFT ((-1))
value DMRES_HIGH ((-4))
value DMRES_LOW ((-2))
value DMRES_MEDIUM ((-3))
value DMTT_BITMAP (1)
value DMTT_DOWNLOAD (2)
value DMTT_DOWNLOAD_OUTLINE (4)
value DMTT_SUBDEV (3)
value DM_BITSPERPEL (0x00040000L)
value DM_COLLATE (0x00008000L)
value DM_COLOR (0x00000800L)
value DM_COPIES (0x00000100L)
value DM_COPY (2)
value DM_DEFAULTSOURCE (0x00000200L)
value DM_DISPLAYFIXEDOUTPUT (0x20000000L)
value DM_DISPLAYFLAGS (0x00200000L)
value DM_DISPLAYFREQUENCY (0x00400000L)
value DM_DISPLAYORIENTATION (0x00000080L)
value DM_DITHERTYPE (0x04000000L)
value DM_DUPLEX (0x00001000L)
value DM_FORMNAME (0x00010000L)
value DM_GETDEFID ((WM_USER+0))
value DM_ICMINTENT (0x01000000L)
value DM_ICMMETHOD (0x00800000L)
value DM_INTERLACED (0x00000002)
value DM_IN_BUFFER (DM_MODIFY)
value DM_IN_PROMPT (DM_PROMPT)
value DM_LOGPIXELS (0x00020000L)
value DM_MEDIATYPE (0x02000000L)
value DM_MODIFY (8)
value DM_NUP (0x00000040L)
value DM_ORIENTATION (0x00000001L)
value DM_OUT_BUFFER (DM_COPY)
value DM_OUT_DEFAULT (DM_UPDATE)
value DM_PANNINGHEIGHT (0x10000000L)
value DM_PANNINGWIDTH (0x08000000L)
value DM_PAPERLENGTH (0x00000004L)
value DM_PAPERSIZE (0x00000002L)
value DM_PAPERWIDTH (0x00000008L)
value DM_PELSHEIGHT (0x00100000L)
value DM_PELSWIDTH (0x00080000L)
value DM_POINTERHITTEST (0x0250)
value DM_POSITION (0x00000020L)
value DM_PRINTQUALITY (0x00000400L)
value DM_PROMPT (4)
value DM_REPOSITION ((WM_USER+2))
value DM_SCALE (0x00000010L)
value DM_SETDEFID ((WM_USER+1))
value DM_SPECVERSION (0x0401)
value DM_TTOPTION (0x00004000L)
value DM_UPDATE (1)
value DM_YRESOLUTION (0x00002000L)
value DNS_ERROR_ADDRESS_REQUIRED (9573)
value DNS_ERROR_ALIAS_LOOP (9722)
value DNS_ERROR_AUTOZONE_ALREADY_EXISTS (9610)
value DNS_ERROR_AXFR (9752)
value DNS_ERROR_BACKGROUND_LOADING (9568)
value DNS_ERROR_BAD_KEYMASTER (9122)
value DNS_ERROR_BAD_PACKET (9502)
value DNS_ERROR_CANNOT_FIND_ROOT_HINTS (9564)
value DNS_ERROR_CLIENT_SUBNET_ALREADY_EXISTS (9977)
value DNS_ERROR_CLIENT_SUBNET_DOES_NOT_EXIST (9976)
value DNS_ERROR_CLIENT_SUBNET_IS_ACCESSED (9975)
value DNS_ERROR_CNAME_COLLISION (9709)
value DNS_ERROR_CNAME_LOOP (9707)
value DNS_ERROR_DATABASE_BASE (9700)
value DNS_ERROR_DATAFILE_BASE (9650)
value DNS_ERROR_DATAFILE_OPEN_FAILURE (9653)
value DNS_ERROR_DATAFILE_PARSING (9655)
value DNS_ERROR_DEFAULT_SCOPE (9960)
value DNS_ERROR_DEFAULT_VIRTUALIZATION_INSTANCE (9925)
value DNS_ERROR_DEFAULT_ZONESCOPE (9953)
value DNS_ERROR_DELEGATION_REQUIRED (9571)
value DNS_ERROR_DNAME_COLLISION (9721)
value DNS_ERROR_DNSSEC_BASE (9100)
value DNS_ERROR_DNSSEC_IS_DISABLED (9125)
value DNS_ERROR_DP_ALREADY_ENLISTED (9904)
value DNS_ERROR_DP_ALREADY_EXISTS (9902)
value DNS_ERROR_DP_BASE (9900)
value DNS_ERROR_DP_DOES_NOT_EXIST (9901)
value DNS_ERROR_DP_FSMO_ERROR (9906)
value DNS_ERROR_DP_NOT_AVAILABLE (9905)
value DNS_ERROR_DP_NOT_ENLISTED (9903)
value DNS_ERROR_DS_UNAVAILABLE (9717)
value DNS_ERROR_DS_ZONE_ALREADY_EXISTS (9718)
value DNS_ERROR_DWORD_VALUE_TOO_LARGE (9567)
value DNS_ERROR_DWORD_VALUE_TOO_SMALL (9566)
value DNS_ERROR_FILE_WRITEBACK_FAILED (9654)
value DNS_ERROR_FORWARDER_ALREADY_EXISTS (9619)
value DNS_ERROR_GENERAL_API_BASE (9550)
value DNS_ERROR_INCONSISTENT_ROOT_HINTS (9565)
value DNS_ERROR_INVAILD_VIRTUALIZATION_INSTANCE_NAME (9924)
value DNS_ERROR_INVALID_CLIENT_SUBNET_NAME (9984)
value DNS_ERROR_INVALID_DATA (ERROR_INVALID_DATA)
value DNS_ERROR_INVALID_DATAFILE_NAME (9652)
value DNS_ERROR_INVALID_INITIAL_ROLLOVER_OFFSET (9115)
value DNS_ERROR_INVALID_IP_ADDRESS (9552)
value DNS_ERROR_INVALID_KEY_SIZE (9106)
value DNS_ERROR_INVALID_NAME (ERROR_INVALID_NAME)
value DNS_ERROR_INVALID_NAME_CHAR (9560)
value DNS_ERROR_INVALID_POLICY_TABLE (9572)
value DNS_ERROR_INVALID_PROPERTY (9553)
value DNS_ERROR_INVALID_ROLLOVER_PERIOD (9114)
value DNS_ERROR_INVALID_SCOPE_NAME (9958)
value DNS_ERROR_INVALID_SCOPE_OPERATION (9961)
value DNS_ERROR_INVALID_SIGNATURE_VALIDITY_PERIOD (9123)
value DNS_ERROR_INVALID_TYPE (9551)
value DNS_ERROR_INVALID_XML (9126)
value DNS_ERROR_INVALID_ZONESCOPE_NAME (9954)
value DNS_ERROR_INVALID_ZONE_OPERATION (9603)
value DNS_ERROR_INVALID_ZONE_TYPE (9611)
value DNS_ERROR_KEYMASTER_REQUIRED (9101)
value DNS_ERROR_KSP_DOES_NOT_SUPPORT_PROTECTION (9108)
value DNS_ERROR_KSP_NOT_ACCESSIBLE (9112)
value DNS_ERROR_LOAD_ZONESCOPE_FAILED (9956)
value DNS_ERROR_MASK (0x00002328)
value DNS_ERROR_NAME_DOES_NOT_EXIST (9714)
value DNS_ERROR_NAME_NOT_IN_ZONE (9706)
value DNS_ERROR_NBSTAT_INIT_FAILED (9617)
value DNS_ERROR_NEED_SECONDARY_ADDRESSES (9614)
value DNS_ERROR_NEED_WINS_SERVERS (9616)
value DNS_ERROR_NODE_CREATION_FAILED (9703)
value DNS_ERROR_NODE_IS_CNAME (9708)
value DNS_ERROR_NODE_IS_DNAME (9720)
value DNS_ERROR_NON_RFC_NAME (9556)
value DNS_ERROR_NOT_ALLOWED_ON_ACTIVE_SKD (9119)
value DNS_ERROR_NOT_ALLOWED_ON_RODC (9569)
value DNS_ERROR_NOT_ALLOWED_ON_ROOT_SERVER (9562)
value DNS_ERROR_NOT_ALLOWED_ON_SIGNED_ZONE (9102)
value DNS_ERROR_NOT_ALLOWED_ON_UNSIGNED_ZONE (9121)
value DNS_ERROR_NOT_ALLOWED_ON_ZSK (9118)
value DNS_ERROR_NOT_ALLOWED_UNDER_DELEGATION (9563)
value DNS_ERROR_NOT_ALLOWED_UNDER_DNAME (9570)
value DNS_ERROR_NOT_ALLOWED_WITH_ZONESCOPES (9955)
value DNS_ERROR_NOT_ENOUGH_SIGNING_KEY_DESCRIPTORS (9104)
value DNS_ERROR_NOT_UNIQUE (9555)
value DNS_ERROR_NO_BOOTFILE_IF_DS_ZONE (9719)
value DNS_ERROR_NO_CREATE_CACHE_DATA (9713)
value DNS_ERROR_NO_DNS_SERVERS (9852)
value DNS_ERROR_NO_MEMORY (ERROR_OUTOFMEMORY)
value DNS_ERROR_NO_PACKET (9503)
value DNS_ERROR_NO_TCPIP (9851)
value DNS_ERROR_NO_VALID_TRUST_ANCHORS (9127)
value DNS_ERROR_NO_ZONE_INFO (9602)
value DNS_ERROR_NUMERIC_NAME (9561)
value DNS_ERROR_OPERATION_BASE (9750)
value DNS_ERROR_PACKET_FMT_BASE (9500)
value DNS_ERROR_POLICY_ALREADY_EXISTS (9971)
value DNS_ERROR_POLICY_DOES_NOT_EXIST (9972)
value DNS_ERROR_POLICY_INVALID_CRITERIA (9973)
value DNS_ERROR_POLICY_INVALID_CRITERIA_CLIENT_SUBNET (9990)
value DNS_ERROR_POLICY_INVALID_CRITERIA_FQDN (9994)
value DNS_ERROR_POLICY_INVALID_CRITERIA_INTERFACE (9993)
value DNS_ERROR_POLICY_INVALID_CRITERIA_NETWORK_PROTOCOL (9992)
value DNS_ERROR_POLICY_INVALID_CRITERIA_QUERY_TYPE (9995)
value DNS_ERROR_POLICY_INVALID_CRITERIA_TIME_OF_DAY (9996)
value DNS_ERROR_POLICY_INVALID_CRITERIA_TRANSPORT_PROTOCOL (9991)
value DNS_ERROR_POLICY_INVALID_NAME (9982)
value DNS_ERROR_POLICY_INVALID_SETTINGS (9974)
value DNS_ERROR_POLICY_INVALID_WEIGHT (9981)
value DNS_ERROR_POLICY_LOCKED (9980)
value DNS_ERROR_POLICY_MISSING_CRITERIA (9983)
value DNS_ERROR_POLICY_PROCESSING_ORDER_INVALID (9985)
value DNS_ERROR_POLICY_SCOPE_MISSING (9986)
value DNS_ERROR_POLICY_SCOPE_NOT_ALLOWED (9987)
value DNS_ERROR_PRIMARY_REQUIRES_DATAFILE (9651)
value DNS_ERROR_RCODE (9504)
value DNS_ERROR_RCODE_BADKEY (9017)
value DNS_ERROR_RCODE_BADSIG (9016)
value DNS_ERROR_RCODE_BADTIME (9018)
value DNS_ERROR_RCODE_FORMAT_ERROR (9001)
value DNS_ERROR_RCODE_LAST (DNS_ERROR_RCODE_BADTIME)
value DNS_ERROR_RCODE_NAME_ERROR (9003)
value DNS_ERROR_RCODE_NOTAUTH (9009)
value DNS_ERROR_RCODE_NOTZONE (9010)
value DNS_ERROR_RCODE_NOT_IMPLEMENTED (9004)
value DNS_ERROR_RCODE_NO_ERROR (NO_ERROR)
value DNS_ERROR_RCODE_NXRRSET (9008)
value DNS_ERROR_RCODE_REFUSED (9005)
value DNS_ERROR_RCODE_SERVER_FAILURE (9002)
value DNS_ERROR_RCODE_YXDOMAIN (9006)
value DNS_ERROR_RCODE_YXRRSET (9007)
value DNS_ERROR_RECORD_ALREADY_EXISTS (9711)
value DNS_ERROR_RECORD_DOES_NOT_EXIST (9701)
value DNS_ERROR_RECORD_FORMAT (9702)
value DNS_ERROR_RECORD_ONLY_AT_ZONE_ROOT (9710)
value DNS_ERROR_RECORD_TIMED_OUT (9705)
value DNS_ERROR_RESPONSE_CODES_BASE (9000)
value DNS_ERROR_ROLLOVER_ALREADY_QUEUED (9120)
value DNS_ERROR_ROLLOVER_IN_PROGRESS (9116)
value DNS_ERROR_ROLLOVER_NOT_POKEABLE (9128)
value DNS_ERROR_RRL_INVALID_LEAK_RATE (9916)
value DNS_ERROR_RRL_INVALID_TC_RATE (9915)
value DNS_ERROR_RRL_INVALID_WINDOW_SIZE (9912)
value DNS_ERROR_RRL_LEAK_RATE_LESSTHAN_TC_RATE (9917)
value DNS_ERROR_RRL_NOT_ENABLED (9911)
value DNS_ERROR_SCOPE_ALREADY_EXISTS (9963)
value DNS_ERROR_SCOPE_DOES_NOT_EXIST (9959)
value DNS_ERROR_SCOPE_LOCKED (9962)
value DNS_ERROR_SECONDARY_DATA (9712)
value DNS_ERROR_SECONDARY_REQUIRES_MASTER_IP (9612)
value DNS_ERROR_SECURE_BASE (9800)
value DNS_ERROR_SERVERSCOPE_IS_REFERENCED (9988)
value DNS_ERROR_SETUP_BASE (9850)
value DNS_ERROR_SIGNING_KEY_NOT_ACCESSIBLE (9107)
value DNS_ERROR_SOA_DELETE_INVALID (9618)
value DNS_ERROR_STANDBY_KEY_NOT_PRESENT (9117)
value DNS_ERROR_SUBNET_ALREADY_EXISTS (9979)
value DNS_ERROR_SUBNET_DOES_NOT_EXIST (9978)
value DNS_ERROR_TOO_MANY_SKDS (9113)
value DNS_ERROR_TRY_AGAIN_LATER (9554)
value DNS_ERROR_UNEXPECTED_CNG_ERROR (9110)
value DNS_ERROR_UNEXPECTED_DATA_PROTECTION_ERROR (9109)
value DNS_ERROR_UNKNOWN_RECORD_TYPE (9704)
value DNS_ERROR_UNKNOWN_SIGNING_PARAMETER_VERSION (9111)
value DNS_ERROR_UNSECURE_PACKET (9505)
value DNS_ERROR_UNSUPPORTED_ALGORITHM (9105)
value DNS_ERROR_VIRTUALIZATION_INSTANCE_ALREADY_EXISTS (9921)
value DNS_ERROR_VIRTUALIZATION_INSTANCE_DOES_NOT_EXIST (9922)
value DNS_ERROR_VIRTUALIZATION_TREE_LOCKED (9923)
value DNS_ERROR_WINS_INIT_FAILED (9615)
value DNS_ERROR_ZONESCOPE_ALREADY_EXISTS (9951)
value DNS_ERROR_ZONESCOPE_DOES_NOT_EXIST (9952)
value DNS_ERROR_ZONESCOPE_FILE_WRITEBACK_FAILED (9957)
value DNS_ERROR_ZONESCOPE_IS_REFERENCED (9989)
value DNS_ERROR_ZONE_ALREADY_EXISTS (9609)
value DNS_ERROR_ZONE_BASE (9600)
value DNS_ERROR_ZONE_CONFIGURATION_ERROR (9604)
value DNS_ERROR_ZONE_CREATION_FAILED (9608)
value DNS_ERROR_ZONE_DOES_NOT_EXIST (9601)
value DNS_ERROR_ZONE_HAS_NO_NS_RECORDS (9606)
value DNS_ERROR_ZONE_HAS_NO_SOA_RECORD (9605)
value DNS_ERROR_ZONE_IS_SHUTDOWN (9621)
value DNS_ERROR_ZONE_LOCKED (9607)
value DNS_ERROR_ZONE_LOCKED_FOR_SIGNING (9622)
value DNS_ERROR_ZONE_NOT_SECONDARY (9613)
value DNS_ERROR_ZONE_REQUIRES_MASTER_IP (9620)
value DNS_FILTEROFF (0x0008)
value DNS_FILTERON (0x0004)
value DNS_INFO_ADDED_LOCAL_WINS (9753)
value DNS_INFO_AXFR_COMPLETE (9751)
value DNS_INFO_NO_RECORDS (9501)
value DNS_REGISTER (0x0001)
value DNS_REQUEST_PENDING (9506)
value DNS_STATUS_CONTINUE_NEEDED (9801)
value DNS_STATUS_DOTTED_NAME (9558)
value DNS_STATUS_FQDN (9557)
value DNS_STATUS_PACKET_UNSECURE (DNS_ERROR_UNSECURE_PACKET)
value DNS_STATUS_SINGLE_PART_NAME (9559)
value DNS_UNREGISTER (0x0002)
value DNS_WARNING_DOMAIN_UNDELETED (9716)
value DNS_WARNING_PTR_CREATE_FAILED (9715)
value DN_DEFAULTPRN (0x0001)
value DOCKINFO_DOCKED ((0x2))
value DOCKINFO_UNDOCKED ((0x1))
value DOCKINFO_USER_DOCKED ((DOCKINFO_USER_SUPPLIED | DOCKINFO_DOCKED))
value DOCKINFO_USER_SUPPLIED ((0x4))
value DOCKINFO_USER_UNDOCKED ((DOCKINFO_USER_SUPPLIED | DOCKINFO_UNDOCKED))
value DOF_DIRECTORY (0x8003)
value DOF_DOCUMENT (0x8002)
value DOF_EXECUTABLE (0x8001)
value DOF_MULTIPLE (0x8004)
value DOF_PROGMAN (0x0001)
value DOF_SHELLDATA (0x0002)
value DOMAIN_ALIAS_RID_ACCESS_CONTROL_ASSISTANCE_OPS ((0x00000243L))
value DOMAIN_ALIAS_RID_ACCOUNT_OPS ((0x00000224L))
value DOMAIN_ALIAS_RID_ADMINS ((0x00000220L))
value DOMAIN_ALIAS_RID_AUTHORIZATIONACCESS ((0x00000230L))
value DOMAIN_ALIAS_RID_BACKUP_OPS ((0x00000227L))
value DOMAIN_ALIAS_RID_CACHEABLE_PRINCIPALS_GROUP ((0x0000023BL))
value DOMAIN_ALIAS_RID_CERTSVC_DCOM_ACCESS_GROUP ((0x0000023EL))
value DOMAIN_ALIAS_RID_CRYPTO_OPERATORS ((0x00000239L))
value DOMAIN_ALIAS_RID_DCOM_USERS ((0x00000232L))
value DOMAIN_ALIAS_RID_DEFAULT_ACCOUNT ((0x00000245L))
value DOMAIN_ALIAS_RID_DEVICE_OWNERS ((0x00000247L))
value DOMAIN_ALIAS_RID_EVENT_LOG_READERS_GROUP ((0x0000023DL))
value DOMAIN_ALIAS_RID_GUESTS ((0x00000222L))
value DOMAIN_ALIAS_RID_HYPER_V_ADMINS ((0x00000242L))
value DOMAIN_ALIAS_RID_INCOMING_FOREST_TRUST_BUILDERS ((0x0000022DL))
value DOMAIN_ALIAS_RID_IUSERS ((0x00000238L))
value DOMAIN_ALIAS_RID_LOGGING_USERS ((0x0000022FL))
value DOMAIN_ALIAS_RID_MONITORING_USERS ((0x0000022EL))
value DOMAIN_ALIAS_RID_NETWORK_CONFIGURATION_OPS ((0x0000022CL))
value DOMAIN_ALIAS_RID_NON_CACHEABLE_PRINCIPALS_GROUP ((0x0000023CL))
value DOMAIN_ALIAS_RID_POWER_USERS ((0x00000223L))
value DOMAIN_ALIAS_RID_PRINT_OPS ((0x00000226L))
value DOMAIN_ALIAS_RID_RAS_SERVERS ((0x00000229L))
value DOMAIN_ALIAS_RID_RDS_ENDPOINT_SERVERS ((0x00000240L))
value DOMAIN_ALIAS_RID_RDS_MANAGEMENT_SERVERS ((0x00000241L))
value DOMAIN_ALIAS_RID_RDS_REMOTE_ACCESS_SERVERS ((0x0000023FL))
value DOMAIN_ALIAS_RID_REMOTE_DESKTOP_USERS ((0x0000022BL))
value DOMAIN_ALIAS_RID_REMOTE_MANAGEMENT_USERS ((0x00000244L))
value DOMAIN_ALIAS_RID_REPLICATOR ((0x00000228L))
value DOMAIN_ALIAS_RID_STORAGE_REPLICA_ADMINS ((0x00000246L))
value DOMAIN_ALIAS_RID_SYSTEM_OPS ((0x00000225L))
value DOMAIN_ALIAS_RID_TS_LICENSE_SERVERS ((0x00000231L))
value DOMAIN_ALIAS_RID_USERS ((0x00000221L))
value DOMAIN_GROUP_RID_ADMINS ((0x00000200L))
value DOMAIN_GROUP_RID_AUTHORIZATION_DATA_CONTAINS_CLAIMS ((0x000001F1L))
value DOMAIN_GROUP_RID_AUTHORIZATION_DATA_IS_COMPOUNDED ((0x000001F0L))
value DOMAIN_GROUP_RID_CDC_RESERVED ((0x0000020CL))
value DOMAIN_GROUP_RID_CERT_ADMINS ((0x00000205L))
value DOMAIN_GROUP_RID_CLONEABLE_CONTROLLERS ((0x0000020AL))
value DOMAIN_GROUP_RID_COMPUTERS ((0x00000203L))
value DOMAIN_GROUP_RID_CONTROLLERS ((0x00000204L))
value DOMAIN_GROUP_RID_ENTERPRISE_ADMINS ((0x00000207L))
value DOMAIN_GROUP_RID_ENTERPRISE_KEY_ADMINS ((0x0000020FL))
value DOMAIN_GROUP_RID_ENTERPRISE_READONLY_DOMAIN_CONTROLLERS ((0x000001F2L))
value DOMAIN_GROUP_RID_GUESTS ((0x00000202L))
value DOMAIN_GROUP_RID_KEY_ADMINS ((0x0000020EL))
value DOMAIN_GROUP_RID_POLICY_ADMINS ((0x00000208L))
value DOMAIN_GROUP_RID_PROTECTED_USERS ((0x0000020DL))
value DOMAIN_GROUP_RID_READONLY_CONTROLLERS ((0x00000209L))
value DOMAIN_GROUP_RID_SCHEMA_ADMINS ((0x00000206L))
value DOMAIN_GROUP_RID_USERS ((0x00000201L))
value DOMAIN_USER_RID_ADMIN ((0x000001F4L))
value DOMAIN_USER_RID_DEFAULT_ACCOUNT ((0x000001F7L))
value DOMAIN_USER_RID_GUEST ((0x000001F5L))
value DOMAIN_USER_RID_KRBTGT ((0x000001F6L))
value DOMAIN_USER_RID_MAX ((0x000003E7L))
value DOMAIN_USER_RID_WDAG_ACCOUNT ((0x000001F8L))
value DONT_RESOLVE_DLL_REFERENCES (0x00000001)
value DOUBLE_CLICK (0x0002)
value DOWNLOADFACE (514)
value DOWNLOADHEADER (4111)
value DO_DROPFILE (0x454C4946L)
value DO_PRINTFILE (0x544E5250L)
value DPD_DELETE_ALL_FILES (0x00000004)
value DPD_DELETE_SPECIFIC_VERSION (0x00000002)
value DPD_DELETE_UNUSED_FILES (0x00000001)
value DPI_AWARENESS_CONTEXT_PER_MONITOR_AWARE (((DPI_AWARENESS_CONTEXT)-3))
value DPI_AWARENESS_CONTEXT_SYSTEM_AWARE (((DPI_AWARENESS_CONTEXT)-2))
value DPI_AWARENESS_CONTEXT_UNAWARE (((DPI_AWARENESS_CONTEXT)-1))
value DPI_AWARENESS_CONTEXT_UNAWARE_GDISCALED (((DPI_AWARENESS_CONTEXT)-5))
value DRAFTMODE (7)
value DRAFT_QUALITY (1)
value DRAGDROP_E_ALREADYREGISTERED (_HRESULT_TYPEDEF_(0x80040101L))
value DRAGDROP_E_CONCURRENT_DRAG_ATTEMPTED (_HRESULT_TYPEDEF_(0x80040103L))
value DRAGDROP_E_FIRST (0x80040100L)
value DRAGDROP_E_INVALIDHWND (_HRESULT_TYPEDEF_(0x80040102L))
value DRAGDROP_E_LAST (0x8004010FL)
value DRAGDROP_E_NOTREGISTERED (_HRESULT_TYPEDEF_(0x80040100L))
value DRAGDROP_S_CANCEL (_HRESULT_TYPEDEF_(0x00040101L))
value DRAGDROP_S_DROP (_HRESULT_TYPEDEF_(0x00040100L))
value DRAGDROP_S_FIRST (0x00040100L)
value DRAGDROP_S_LAST (0x0004010FL)
value DRAGDROP_S_USEDEFAULTCURSORS (_HRESULT_TYPEDEF_(0x00040102L))
value DRAWPATTERNRECT (25)
value DRIVERVERSION (0)
value DRIVER_KERNELMODE (0x00000001)
value DRIVER_USERMODE (0x00000002)
value DRIVE_CDROM (5)
value DRIVE_FIXED (3)
value DRIVE_NO_ROOT_DIR (1)
value DRIVE_RAMDISK (6)
value DRIVE_REMOTE (4)
value DRIVE_REMOVABLE (2)
value DRIVE_UNKNOWN (0)
value DROPEFFECT_COPY (( 1 ))
value DROPEFFECT_LINK (( 4 ))
value DROPEFFECT_MOVE (( 2 ))
value DROPEFFECT_NONE (( 0 ))
value DROPEFFECT_SCROLL (( 0x80000000 ))
value DRVCNF_CANCEL (0x0000)
value DRVCNF_OK (0x0001)
value DRVCNF_RESTART (0x0002)
value DRV_CANCEL (DRVCNF_CANCEL)
value DRV_CLOSE (0x0004)
value DRV_CONFIGURE (0x0007)
value DRV_DISABLE (0x0005)
value DRV_ENABLE (0x0002)
value DRV_EXITSESSION (0x000B)
value DRV_FREE (0x0006)
value DRV_INSTALL (0x0009)
value DRV_LOAD (0x0001)
value DRV_MCI_FIRST (DRV_RESERVED)
value DRV_MCI_LAST ((DRV_RESERVED + 0xFFF))
value DRV_OK (DRVCNF_OK)
value DRV_OPEN (0x0003)
value DRV_POWER (0x000F)
value DRV_QUERYCONFIGURE (0x0008)
value DRV_REMOVE (0x000A)
value DRV_RESERVED (0x0800)
value DRV_RESTART (DRVCNF_RESTART)
value DRV_USER (0x4000)
value DSPRINT_PENDING (0x80000000)
value DSPRINT_PUBLISH (0x00000001)
value DSPRINT_REPUBLISH (0x00000008)
value DSPRINT_UNPUBLISH (0x00000004)
value DSPRINT_UPDATE (0x00000002)
value DSS_DISABLED (0x0020)
value DSS_HIDEPREFIX (0x0200)
value DSS_MONO (0x0080)
value DSS_NORMAL (0x0000)
value DSS_PREFIXONLY (0x0400)
value DSS_RIGHT (0x8000)
value DSS_UNION (0x0010)
value DSTINVERT ((DWORD)0x00550009)
value DST_BITMAP (0x0004)
value DST_COMPLEX (0x0000)
value DST_ICON (0x0003)
value DST_PREFIXTEXT (0x0002)
value DST_TEXT (0x0001)
value DS_ABSALIGN (0x01L)
value DS_CENTER (0x0800L)
value DS_CENTERMOUSE (0x1000L)
value DS_CONTEXTHELP (0x2000L)
value DS_CONTROL (0x0400L)
value DS_FIXEDSYS (0x0008L)
value DS_LOCALEDIT (0x20L)
value DS_MODALFRAME (0x80L)
value DS_NOFAILCREATE (0x0010L)
value DS_NOIDLEMSG (0x100L)
value DS_SETFONT (0x40L)
value DS_SETFOREGROUND (0x200L)
value DS_SHELLFONT ((DS_SETFONT | DS_FIXEDSYS))
value DS_SYSMODAL (0x02L)
value DS_S_SUCCESS (NO_ERROR)
value DTR_CONTROL_DISABLE (0x00)
value DTR_CONTROL_ENABLE (0x01)
value DTR_CONTROL_HANDSHAKE (0x02)
value DT_BOTTOM (0x00000008)
value DT_CALCRECT (0x00000400)
value DT_CENTER (0x00000001)
value DT_CHARSTREAM (4)
value DT_DISPFILE (6)
value DT_EDITCONTROL (0x00002000)
value DT_END_ELLIPSIS (0x00008000)
value DT_EXPANDTABS (0x00000040)
value DT_EXTERNALLEADING (0x00000200)
value DT_HIDEPREFIX (0x00100000)
value DT_INTERNAL (0x00001000)
value DT_LEFT (0x00000000)
value DT_METAFILE (5)
value DT_MODIFYSTRING (0x00010000)
value DT_NOCLIP (0x00000100)
value DT_NOFULLWIDTHCHARBREAK (0x00080000)
value DT_NOPREFIX (0x00000800)
value DT_PATH_ELLIPSIS (0x00004000)
value DT_PLOTTER (0)
value DT_PREFIXONLY (0x00200000)
value DT_RASCAMERA (3)
value DT_RASDISPLAY (1)
value DT_RASPRINTER (2)
value DT_RIGHT (0x00000002)
value DT_RTLREADING (0x00020000)
value DT_SINGLELINE (0x00000020)
value DT_TABSTOP (0x00000080)
value DT_TOP (0x00000000)
value DT_VCENTER (0x00000004)
value DT_WORDBREAK (0x00000010)
value DT_WORD_ELLIPSIS (0x00040000)
value DUPLICATE (0x06)
value DUPLICATE_CLOSE_SOURCE (0x00000001)
value DUPLICATE_DEREG (0x07)
value DUPLICATE_EXTENTS_DATA_EX_ASYNC (0x00000002)
value DUPLICATE_EXTENTS_DATA_EX_SOURCE_ATOMIC (0x00000001)
value DUPLICATE_SAME_ACCESS (0x00000002)
value DV_E_CLIPFORMAT (_HRESULT_TYPEDEF_(0x8004006AL))
value DV_E_DVASPECT (_HRESULT_TYPEDEF_(0x8004006BL))
value DV_E_DVTARGETDEVICE (_HRESULT_TYPEDEF_(0x80040065L))
value DV_E_DVTARGETDEVICE_SIZE (_HRESULT_TYPEDEF_(0x8004006CL))
value DV_E_FORMATETC (_HRESULT_TYPEDEF_(0x80040064L))
value DV_E_LINDEX (_HRESULT_TYPEDEF_(0x80040068L))
value DV_E_NOIVIEWOBJECT (_HRESULT_TYPEDEF_(0x8004006DL))
value DV_E_STATDATA (_HRESULT_TYPEDEF_(0x80040067L))
value DV_E_STGMEDIUM (_HRESULT_TYPEDEF_(0x80040066L))
value DV_E_TYMED (_HRESULT_TYPEDEF_(0x80040069L))
value DWLP_MSGRESULT (0)
value DWMERR_CATASTROPHIC_FAILURE (_HRESULT_TYPEDEF_(0x88980702L))
value DWMERR_STATE_TRANSITION_FAILED (_HRESULT_TYPEDEF_(0x88980700L))
value DWMERR_THEME_FAILED (_HRESULT_TYPEDEF_(0x88980701L))
value DWM_E_ADAPTER_NOT_FOUND (_HRESULT_TYPEDEF_(0x80263005L))
value DWM_E_COMPOSITIONDISABLED (_HRESULT_TYPEDEF_(0x80263001L))
value DWM_E_NOT_QUEUING_PRESENTS (_HRESULT_TYPEDEF_(0x80263004L))
value DWM_E_NO_REDIRECTION_SURFACE_AVAILABLE (_HRESULT_TYPEDEF_(0x80263003L))
value DWM_E_REMOTING_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80263002L))
value DWM_E_TEXTURE_TOO_LARGE (_HRESULT_TYPEDEF_(0x80263007L))
value DWM_S_GDI_REDIRECTION_SURFACE (_HRESULT_TYPEDEF_(0x00263005L))
value DWM_S_GDI_REDIRECTION_SURFACE_BLT_VIA_GDI (_HRESULT_TYPEDEF_(0x00263008L))
value DWRITE_E_ALREADYREGISTERED (_HRESULT_TYPEDEF_(0x88985006L))
value DWRITE_E_CACHEFORMAT (_HRESULT_TYPEDEF_(0x88985007L))
value DWRITE_E_CACHEVERSION (_HRESULT_TYPEDEF_(0x88985008L))
value DWRITE_E_DOWNLOADCANCELLED (_HRESULT_TYPEDEF_(0x8898500EL))
value DWRITE_E_DOWNLOADFAILED (_HRESULT_TYPEDEF_(0x8898500FL))
value DWRITE_E_FILEACCESS (_HRESULT_TYPEDEF_(0x88985004L))
value DWRITE_E_FILEFORMAT (_HRESULT_TYPEDEF_(0x88985000L))
value DWRITE_E_FILENOTFOUND (_HRESULT_TYPEDEF_(0x88985003L))
value DWRITE_E_FLOWDIRECTIONCONFLICTS (_HRESULT_TYPEDEF_(0x8898500BL))
value DWRITE_E_FONTCOLLECTIONOBSOLETE (_HRESULT_TYPEDEF_(0x88985005L))
value DWRITE_E_NOCOLOR (_HRESULT_TYPEDEF_(0x8898500CL))
value DWRITE_E_NOFONT (_HRESULT_TYPEDEF_(0x88985002L))
value DWRITE_E_REMOTEFONT (_HRESULT_TYPEDEF_(0x8898500DL))
value DWRITE_E_TEXTRENDERERINCOMPATIBLE (_HRESULT_TYPEDEF_(0x8898500AL))
value DWRITE_E_TOOMANYDOWNLOADS (_HRESULT_TYPEDEF_(0x88985010L))
value DWRITE_E_UNEXPECTED (_HRESULT_TYPEDEF_(0x88985001L))
value DWRITE_E_UNSUPPORTEDOPERATION (_HRESULT_TYPEDEF_(0x88985009L))
value DXCORE_ERROR_EVENT_NOT_UNREGISTERED (_HRESULT_TYPEDEF_(0x88800001L))
value DXGI_DDI_ERR_NONEXCLUSIVE (_HRESULT_TYPEDEF_(0x887B0003L))
value DXGI_DDI_ERR_UNSUPPORTED (_HRESULT_TYPEDEF_(0x887B0002L))
value DXGI_DDI_ERR_WASSTILLDRAWING (_HRESULT_TYPEDEF_(0x887B0001L))
value DXGI_ERROR_ACCESS_DENIED (_HRESULT_TYPEDEF_(0x887A002BL))
value DXGI_ERROR_ACCESS_LOST (_HRESULT_TYPEDEF_(0x887A0026L))
value DXGI_ERROR_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x887A0036L))
value DXGI_ERROR_CACHE_CORRUPT (_HRESULT_TYPEDEF_(0x887A0033L))
value DXGI_ERROR_CACHE_FULL (_HRESULT_TYPEDEF_(0x887A0034L))
value DXGI_ERROR_CACHE_HASH_COLLISION (_HRESULT_TYPEDEF_(0x887A0035L))
value DXGI_ERROR_CANNOT_PROTECT_CONTENT (_HRESULT_TYPEDEF_(0x887A002AL))
value DXGI_ERROR_DEVICE_HUNG (_HRESULT_TYPEDEF_(0x887A0006L))
value DXGI_ERROR_DEVICE_REMOVED (_HRESULT_TYPEDEF_(0x887A0005L))
value DXGI_ERROR_DEVICE_RESET (_HRESULT_TYPEDEF_(0x887A0007L))
value DXGI_ERROR_DRIVER_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x887A0020L))
value DXGI_ERROR_DYNAMIC_CODE_POLICY_VIOLATION (_HRESULT_TYPEDEF_(0x887A0031L))
value DXGI_ERROR_FRAME_STATISTICS_DISJOINT (_HRESULT_TYPEDEF_(0x887A000BL))
value DXGI_ERROR_GRAPHICS_VIDPN_SOURCE_IN_USE (_HRESULT_TYPEDEF_(0x887A000CL))
value DXGI_ERROR_HW_PROTECTION_OUTOFMEMORY (_HRESULT_TYPEDEF_(0x887A0030L))
value DXGI_ERROR_INVALID_CALL (_HRESULT_TYPEDEF_(0x887A0001L))
value DXGI_ERROR_MODE_CHANGE_IN_PROGRESS (_HRESULT_TYPEDEF_(0x887A0025L))
value DXGI_ERROR_MORE_DATA (_HRESULT_TYPEDEF_(0x887A0003L))
value DXGI_ERROR_MPO_UNPINNED (_HRESULT_TYPEDEF_(0x887A0064L))
value DXGI_ERROR_NAME_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x887A002CL))
value DXGI_ERROR_NONEXCLUSIVE (_HRESULT_TYPEDEF_(0x887A0021L))
value DXGI_ERROR_NON_COMPOSITED_UI (_HRESULT_TYPEDEF_(0x887A0032L))
value DXGI_ERROR_NOT_CURRENT (_HRESULT_TYPEDEF_(0x887A002EL))
value DXGI_ERROR_NOT_CURRENTLY_AVAILABLE (_HRESULT_TYPEDEF_(0x887A0022L))
value DXGI_ERROR_NOT_FOUND (_HRESULT_TYPEDEF_(0x887A0002L))
value DXGI_ERROR_REMOTE_CLIENT_DISCONNECTED (_HRESULT_TYPEDEF_(0x887A0023L))
value DXGI_ERROR_REMOTE_OUTOFMEMORY (_HRESULT_TYPEDEF_(0x887A0024L))
value DXGI_ERROR_RESTRICT_TO_OUTPUT_STALE (_HRESULT_TYPEDEF_(0x887A0029L))
value DXGI_ERROR_SDK_COMPONENT_MISSING (_HRESULT_TYPEDEF_(0x887A002DL))
value DXGI_ERROR_SESSION_DISCONNECTED (_HRESULT_TYPEDEF_(0x887A0028L))
value DXGI_ERROR_UNSUPPORTED (_HRESULT_TYPEDEF_(0x887A0004L))
value DXGI_ERROR_WAIT_TIMEOUT (_HRESULT_TYPEDEF_(0x887A0027L))
value DXGI_ERROR_WAS_STILL_DRAWING (_HRESULT_TYPEDEF_(0x887A000AL))
value DXGI_STATUS_CLIPPED (_HRESULT_TYPEDEF_(0x087A0002L))
value DXGI_STATUS_DDA_WAS_STILL_DRAWING (_HRESULT_TYPEDEF_(0x087A000AL))
value DXGI_STATUS_GRAPHICS_VIDPN_SOURCE_IN_USE (_HRESULT_TYPEDEF_(0x087A0006L))
value DXGI_STATUS_MODE_CHANGED (_HRESULT_TYPEDEF_(0x087A0007L))
value DXGI_STATUS_MODE_CHANGE_IN_PROGRESS (_HRESULT_TYPEDEF_(0x087A0008L))
value DXGI_STATUS_NO_DESKTOP_ACCESS (_HRESULT_TYPEDEF_(0x087A0005L))
value DXGI_STATUS_NO_REDIRECTION (_HRESULT_TYPEDEF_(0x087A0004L))
value DXGI_STATUS_OCCLUDED (_HRESULT_TYPEDEF_(0x087A0001L))
value DXGI_STATUS_PRESENT_REQUIRED (_HRESULT_TYPEDEF_(0x087A002FL))
value DXGI_STATUS_UNOCCLUDED (_HRESULT_TYPEDEF_(0x087A0009L))
value DYNAMIC_EH_CONTINUATION_TARGET_ADD ((0x00000001))
value DYNAMIC_EH_CONTINUATION_TARGET_PROCESSED ((0x00000002))
value DYNAMIC_ENFORCED_ADDRESS_RANGE_ADD ((0x00000001))
value DYNAMIC_ENFORCED_ADDRESS_RANGE_PROCESSED ((0x00000002))
value EACCES (13)
value EADDRINUSE (100)
value EADDRNOTAVAIL (101)
value EAFNOSUPPORT (102)
value EAGAIN (11)
value EALREADY (103)
value EASTEUROPE_CHARSET (238)
value EAS_E_ADMINS_CANNOT_CHANGE_PASSWORD (_HRESULT_TYPEDEF_(0x80550008L))
value EAS_E_ADMINS_HAVE_BLANK_PASSWORD (_HRESULT_TYPEDEF_(0x80550007L))
value EAS_E_CONNECTED_ADMINS_NEED_TO_CHANGE_PASSWORD (_HRESULT_TYPEDEF_(0x8055000BL))
value EAS_E_CURRENT_CONNECTED_USER_NEED_TO_CHANGE_PASSWORD (_HRESULT_TYPEDEF_(0x8055000DL))
value EAS_E_CURRENT_USER_HAS_BLANK_PASSWORD (_HRESULT_TYPEDEF_(0x80550004L))
value EAS_E_LOCAL_CONTROLLED_USERS_CANNOT_CHANGE_PASSWORD (_HRESULT_TYPEDEF_(0x80550009L))
value EAS_E_PASSWORD_POLICY_NOT_ENFORCEABLE_FOR_CONNECTED_ADMINS (_HRESULT_TYPEDEF_(0x8055000AL))
value EAS_E_PASSWORD_POLICY_NOT_ENFORCEABLE_FOR_CURRENT_CONNECTED_USER (_HRESULT_TYPEDEF_(0x8055000CL))
value EAS_E_POLICY_COMPLIANT_WITH_ACTIONS (_HRESULT_TYPEDEF_(0x80550002L))
value EAS_E_POLICY_NOT_MANAGED_BY_OS (_HRESULT_TYPEDEF_(0x80550001L))
value EAS_E_REQUESTED_POLICY_NOT_ENFORCEABLE (_HRESULT_TYPEDEF_(0x80550003L))
value EAS_E_REQUESTED_POLICY_PASSWORD_EXPIRATION_INCOMPATIBLE (_HRESULT_TYPEDEF_(0x80550005L))
value EAS_E_USER_CANNOT_CHANGE_PASSWORD (_HRESULT_TYPEDEF_(0x80550006L))
value EBADF (9)
value EBADMSG (104)
value EBUSY (16)
value ECANCELED (105)
value ECC_CMS_SHARED_INFO (((LPCSTR) 77))
value ECHILD (10)
value ECONNABORTED (106)
value ECONNREFUSED (107)
value ECONNRESET (108)
value EC_DISABLE (ST_BLOCKED)
value EC_ENABLEALL (0)
value EC_ENABLEONE (ST_BLOCKNEXT)
value EC_LEFTMARGIN (0x0001)
value EC_QUERYWAITING (2)
value EC_RIGHTMARGIN (0x0002)
value EC_USEFONTINFO (0xffff)
value EDD_GET_DEVICE_INTERFACE_NAME (0x00000001)
value EDEADLK (36)
value EDEADLOCK (EDEADLK)
value EDESTADDRREQ (109)
value EDGE_BUMP ((BDR_RAISEDOUTER | BDR_SUNKENINNER))
value EDGE_ETCHED ((BDR_SUNKENOUTER | BDR_RAISEDINNER))
value EDGE_RAISED ((BDR_RAISEDOUTER | BDR_RAISEDINNER))
value EDGE_SUNKEN ((BDR_SUNKENOUTER | BDR_SUNKENINNER))
value EDOM (33)
value EDS_RAWMODE (0x00000002)
value EDS_ROTATEDMODE (0x00000004)
value EEXIST (17)
value EFAULT (14)
value EFBIG (27)
value EFSRPC_SECURE_ONLY ((8))
value EFS_COMPATIBILITY_VERSION_NCRYPT_PROTECTOR (5)
value EFS_COMPATIBILITY_VERSION_PFILE_PROTECTOR (6)
value EFS_DROP_ALTERNATE_STREAMS ((0x10))
value EFS_EFS_SUBVER_EFS_CERT (1)
value EFS_METADATA_ADD_USER (0x00000001)
value EFS_METADATA_GENERAL_OP (0x00000008)
value EFS_METADATA_REMOVE_USER (0x00000002)
value EFS_METADATA_REPLACE_USER (0x00000004)
value EFS_PFILE_SUBVER_APPX (3)
value EFS_PFILE_SUBVER_RMS (2)
value EFS_SUBVER_UNKNOWN (0)
value EFS_TRACKED_OFFSET_HEADER_FLAG (0x0001)
value EFS_USE_RECOVERY_KEYS ((0x1))
value EHOSTUNREACH (110)
value EIDRM (111)
value EILSEQ (42)
value EIMES_CANCELCOMPSTRINFOCUS (0x0002)
value EIMES_COMPLETECOMPSTRKILLFOCUS (0x0004)
value EIMES_GETCOMPSTRATONCE (0x0001)
value EINPROGRESS (112)
value EINTR (4)
value EINVAL (22)
value EIO (5)
value EISCONN (113)
value EISDIR (21)
value ELEMENT_STATUS_ACCESS (0x00000008)
value ELEMENT_STATUS_AVOLTAG (0x20000000)
value ELEMENT_STATUS_EXCEPT (0x00000004)
value ELEMENT_STATUS_EXENAB (0x00000010)
value ELEMENT_STATUS_FULL (0x00000001)
value ELEMENT_STATUS_ID_VALID (0x00002000)
value ELEMENT_STATUS_IMPEXP (0x00000002)
value ELEMENT_STATUS_INENAB (0x00000020)
value ELEMENT_STATUS_INVERT (0x00400000)
value ELEMENT_STATUS_LUN_VALID (0x00001000)
value ELEMENT_STATUS_NOT_BUS (0x00008000)
value ELEMENT_STATUS_PRODUCT_DATA (0x00000040)
value ELEMENT_STATUS_PVOLTAG (0x10000000)
value ELEMENT_STATUS_SVALID (0x00800000)
value ELF_CULTURE_LATIN (0)
value ELF_VENDOR_SIZE (4)
value ELF_VERSION (0)
value ELOOP (114)
value EMBDHLP_CREATENOW (0x00000000L)
value EMBDHLP_DELAYCREATE (0x00010000L)
value EMBDHLP_INPROC_HANDLER (0x0000L)
value EMBDHLP_INPROC_SERVER (0x0001L)
value EMFILE (24)
value EMLINK (31)
value EMR_ABORTPATH (68)
value EMR_ALPHABLEND (114)
value EMR_ANGLEARC (41)
value EMR_ARC (45)
value EMR_ARCTO (55)
value EMR_BEGINPATH (59)
value EMR_BITBLT (76)
value EMR_CHORD (46)
value EMR_CLOSEFIGURE (61)
value EMR_COLORCORRECTPALETTE (111)
value EMR_COLORMATCHTOTARGETW (121)
value EMR_CREATEBRUSHINDIRECT (39)
value EMR_CREATECOLORSPACE (99)
value EMR_CREATECOLORSPACEW (122)
value EMR_CREATEDIBPATTERNBRUSHPT (94)
value EMR_CREATEMONOBRUSH (93)
value EMR_CREATEPALETTE (49)
value EMR_CREATEPEN (38)
value EMR_DELETECOLORSPACE (101)
value EMR_DELETEOBJECT (40)
value EMR_ELLIPSE (42)
value EMR_ENDPATH (60)
value EMR_EOF (14)
value EMR_EXCLUDECLIPRECT (29)
value EMR_EXTCREATEFONTINDIRECTW (82)
value EMR_EXTCREATEPEN (95)
value EMR_EXTFLOODFILL (53)
value EMR_EXTSELECTCLIPRGN (75)
value EMR_EXTTEXTOUTA (83)
value EMR_EXTTEXTOUTW (84)
value EMR_FILLPATH (62)
value EMR_FILLRGN (71)
value EMR_FLATTENPATH (65)
value EMR_FRAMERGN (72)
value EMR_GDICOMMENT (70)
value EMR_GLSBOUNDEDRECORD (103)
value EMR_GLSRECORD (102)
value EMR_GRADIENTFILL (118)
value EMR_HEADER (1)
value EMR_INTERSECTCLIPRECT (30)
value EMR_INVERTRGN (73)
value EMR_LINETO (54)
value EMR_MASKBLT (78)
value EMR_MAX (122)
value EMR_MIN (1)
value EMR_MODIFYWORLDTRANSFORM (36)
value EMR_MOVETOEX (27)
value EMR_OFFSETCLIPRGN (26)
value EMR_PAINTRGN (74)
value EMR_PIE (47)
value EMR_PIXELFORMAT (104)
value EMR_PLGBLT (79)
value EMR_POLYBEZIER (2)
value EMR_POLYBEZIERTO (5)
value EMR_POLYDRAW (56)
value EMR_POLYGON (3)
value EMR_POLYLINE (4)
value EMR_POLYLINETO (6)
value EMR_POLYPOLYGON (8)
value EMR_POLYPOLYLINE (7)
value EMR_POLYTEXTOUTA (96)
value EMR_POLYTEXTOUTW (97)
value EMR_REALIZEPALETTE (52)
value EMR_RECTANGLE (43)
value EMR_RESIZEPALETTE (51)
value EMR_RESTOREDC (34)
value EMR_ROUNDRECT (44)
value EMR_SAVEDC (33)
value EMR_SCALEVIEWPORTEXTEX (31)
value EMR_SCALEWINDOWEXTEX (32)
value EMR_SELECTCLIPPATH (67)
value EMR_SELECTOBJECT (37)
value EMR_SELECTPALETTE (48)
value EMR_SETARCDIRECTION (57)
value EMR_SETBKCOLOR (25)
value EMR_SETBKMODE (18)
value EMR_SETBRUSHORGEX (13)
value EMR_SETCOLORADJUSTMENT (23)
value EMR_SETCOLORSPACE (100)
value EMR_SETDIBITSTODEVICE (80)
value EMR_SETICMMODE (98)
value EMR_SETICMPROFILEA (112)
value EMR_SETICMPROFILEW (113)
value EMR_SETLAYOUT (115)
value EMR_SETMAPMODE (17)
value EMR_SETMAPPERFLAGS (16)
value EMR_SETMETARGN (28)
value EMR_SETMITERLIMIT (58)
value EMR_SETPALETTEENTRIES (50)
value EMR_SETPIXELV (15)
value EMR_SETPOLYFILLMODE (19)
value EMR_SETSTRETCHBLTMODE (21)
value EMR_SETTEXTALIGN (22)
value EMR_SETTEXTCOLOR (24)
value EMR_SETVIEWPORTEXTEX (11)
value EMR_SETVIEWPORTORGEX (12)
value EMR_SETWINDOWEXTEX (9)
value EMR_SETWINDOWORGEX (10)
value EMR_SETWORLDTRANSFORM (35)
value EMR_STRETCHBLT (77)
value EMR_STRETCHDIBITS (81)
value EMR_STROKEANDFILLPATH (63)
value EMR_STROKEPATH (64)
value EMR_TRANSPARENTBLT (116)
value EMR_WIDENPATH (66)
value EMSGSIZE (115)
value EMSIS_COMPOSITIONSTRING (0x0001)
value EM_CANUNDO (0x00C6)
value EM_CHARFROMPOS (0x00D7)
value EM_EMPTYUNDOBUFFER (0x00CD)
value EM_ENABLEFEATURE (0x00DA)
value EM_FMTLINES (0x00C8)
value EM_GETFIRSTVISIBLELINE (0x00CE)
value EM_GETHANDLE (0x00BD)
value EM_GETIMESTATUS (0x00D9)
value EM_GETLIMITTEXT (0x00D5)
value EM_GETLINE (0x00C4)
value EM_GETLINECOUNT (0x00BA)
value EM_GETMARGINS (0x00D4)
value EM_GETMODIFY (0x00B8)
value EM_GETPASSWORDCHAR (0x00D2)
value EM_GETRECT (0x00B2)
value EM_GETSEL (0x00B0)
value EM_GETTHUMB (0x00BE)
value EM_GETWORDBREAKPROC (0x00D1)
value EM_LIMITTEXT (0x00C5)
value EM_LINEFROMCHAR (0x00C9)
value EM_LINEINDEX (0x00BB)
value EM_LINELENGTH (0x00C1)
value EM_LINESCROLL (0x00B6)
value EM_POSFROMCHAR (0x00D6)
value EM_REPLACESEL (0x00C2)
value EM_SCROLL (0x00B5)
value EM_SCROLLCARET (0x00B7)
value EM_SETHANDLE (0x00BC)
value EM_SETIMESTATUS (0x00D8)
value EM_SETLIMITTEXT (EM_LIMITTEXT)
value EM_SETMARGINS (0x00D3)
value EM_SETMODIFY (0x00B9)
value EM_SETPASSWORDCHAR (0x00CC)
value EM_SETREADONLY (0x00CF)
value EM_SETRECT (0x00B3)
value EM_SETRECTNP (0x00B4)
value EM_SETSEL (0x00B1)
value EM_SETTABSTOPS (0x00CB)
value EM_SETWORDBREAKPROC (0x00D0)
value EM_UNDO (0x00C7)
value ENABLEDUPLEX (28)
value ENABLEPAIRKERNING (769)
value ENABLERELATIVEWIDTHS (768)
value ENABLE_AUTO_POSITION (0x0100)
value ENABLE_DISABLE_AUTOSAVE (0xD2)
value ENABLE_DISABLE_AUTO_OFFLINE (0xDB)
value ENABLE_ECHO_INPUT (0x0004)
value ENABLE_EXTENDED_FLAGS (0x0080)
value ENABLE_INSERT_MODE (0x0020)
value ENABLE_LINE_INPUT (0x0002)
value ENABLE_LVB_GRID_WORLDWIDE (0x0010)
value ENABLE_MOUSE_INPUT (0x0010)
value ENABLE_PROCESSED_INPUT (0x0001)
value ENABLE_PROCESSED_OUTPUT (0x0001)
value ENABLE_QUICK_EDIT_MODE (0x0040)
value ENABLE_SMART (0xD8)
value ENABLE_VIRTUAL_TERMINAL_INPUT (0x0200)
value ENABLE_VIRTUAL_TERMINAL_PROCESSING (0x0004)
value ENABLE_WINDOW_INPUT (0x0008)
value ENABLE_WRAP_AT_EOL_OUTPUT (0x0002)
value ENAMETOOLONG (38)
value ENCAPSULATED_POSTSCRIPT (4116)
value ENCLAVE_LONG_ID_LENGTH (32)
value ENCLAVE_SHORT_ID_LENGTH (16)
value ENCLAVE_TYPE_SGX (0x00000001)
value ENCLAVE_TYPE_VBS (0x00000010)
value ENCLAVE_TYPE_VBS_BASIC (0x00000011)
value ENCLAVE_VBS_FLAG_DEBUG (0x00000001)
value ENCRYPTED_DATA_INFO_SPARSE_FILE (1)
value ENCRYPTION_FORMAT_DEFAULT ((0x01))
value ENDDOC (11)
value ENDSESSION_CLOSEAPP (0x00000001)
value ENDSESSION_CRITICAL (0x40000000)
value ENDSESSION_LOGOFF (0x80000000)
value END_PATH (4098)
value ENETDOWN (116)
value ENETRESET (117)
value ENETUNREACH (118)
value ENFILE (23)
value ENHANCED_KEY (0x0100)
value ENHMETA_SIGNATURE (0x464D4520)
value ENHMETA_STOCK_OBJECT (0x80000000)
value ENLISTMENT_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | ENLISTMENT_GENERIC_READ | ENLISTMENT_GENERIC_WRITE | ENLISTMENT_GENERIC_EXECUTE))
value ENLISTMENT_GENERIC_EXECUTE ((STANDARD_RIGHTS_EXECUTE | ENLISTMENT_RECOVER | ENLISTMENT_SUBORDINATE_RIGHTS | ENLISTMENT_SUPERIOR_RIGHTS))
value ENLISTMENT_GENERIC_READ ((STANDARD_RIGHTS_READ | ENLISTMENT_QUERY_INFORMATION))
value ENLISTMENT_GENERIC_WRITE ((STANDARD_RIGHTS_WRITE | ENLISTMENT_SET_INFORMATION | ENLISTMENT_RECOVER | ENLISTMENT_SUBORDINATE_RIGHTS | ENLISTMENT_SUPERIOR_RIGHTS))
value ENLISTMENT_MAXIMUM_OPTION (0x00000001)
value ENLISTMENT_QUERY_INFORMATION (( 0x0001 ))
value ENLISTMENT_RECOVER (( 0x0004 ))
value ENLISTMENT_SET_INFORMATION (( 0x0002 ))
value ENLISTMENT_SUBORDINATE_RIGHTS (( 0x0008 ))
value ENLISTMENT_SUPERIOR (0x00000001)
value ENLISTMENT_SUPERIOR_RIGHTS (( 0x0010 ))
value ENOBUFS (119)
value ENODATA (120)
value ENODEV (19)
value ENOENT (2)
value ENOEXEC (8)
value ENOLCK (39)
value ENOLINK (121)
value ENOMEM (12)
value ENOMSG (122)
value ENOPROTOOPT (123)
value ENOSPC (28)
value ENOSR (124)
value ENOSTR (125)
value ENOSYS (40)
value ENOTCONN (126)
value ENOTDIR (20)
value ENOTEMPTY (41)
value ENOTRECOVERABLE (127)
value ENOTSOCK (128)
value ENOTSUP (129)
value ENOTTY (25)
value ENUMPAPERBINS (31)
value ENUMPAPERMETRICS (34)
value ENUMRESLANGPROC (ENUMRESLANGPROCA)
value ENUMRESNAMEPROC (ENUMRESNAMEPROCA)
value ENUMRESTYPEPROC (ENUMRESTYPEPROCA)
value ENUM_ALL_CALENDARS (0xffffffff)
value ENUM_CURRENT_SETTINGS (((DWORD)-1))
value ENUM_E_FIRST (0x800401B0L)
value ENUM_E_LAST (0x800401BFL)
value ENUM_REGISTRY_SETTINGS (((DWORD)-2))
value ENUM_S_FIRST (0x000401B0L)
value ENUM_S_LAST (0x000401BFL)
value ENXIO (6)
value EN_AFTER_PASTE (0x0801)
value EN_ALIGN_LTR_EC (0x0700)
value EN_ALIGN_RTL_EC (0x0701)
value EN_BEFORE_PASTE (0x0800)
value EN_CHANGE (0x0300)
value EN_ERRSPACE (0x0500)
value EN_HSCROLL (0x0601)
value EN_KILLFOCUS (0x0200)
value EN_MAXTEXT (0x0501)
value EN_SETFOCUS (0x0100)
value EN_UPDATE (0x0400)
value EN_VSCROLL (0x0602)
value EOF ((-1))
value EOPNOTSUPP (130)
value EOTHER (131)
value EOVERFLOW (132)
value EOWNERDEAD (133)
value EPERM (1)
value EPIPE (32)
value EPROTO (134)
value EPROTONOSUPPORT (135)
value EPROTOTYPE (136)
value EPSPRINTING (33)
value EPS_SIGNATURE (0x46535045)
value EPT_S_CANT_CREATE (1899)
value EPT_S_CANT_PERFORM_OP (1752)
value EPT_S_INVALID_ENTRY (1751)
value EPT_S_NOT_REGISTERED (1753)
value ERANGE (34)
value EROFS (30)
value ERROR (0)
value ERROR_ABANDON_HIBERFILE (787)
value ERROR_ABIOS_ERROR (538)
value ERROR_ACCESS_AUDIT_BY_POLICY (785)
value ERROR_ACCESS_DENIED (5)
value ERROR_ACCESS_DENIED_APPDATA (502)
value ERROR_ACCESS_DISABLED_BY_POLICY (1260)
value ERROR_ACCESS_DISABLED_NO_SAFER_UI_BY_POLICY (786)
value ERROR_ACCESS_DISABLED_WEBBLADE (1277)
value ERROR_ACCESS_DISABLED_WEBBLADE_TAMPER (1278)
value ERROR_ACCOUNT_DISABLED (1331)
value ERROR_ACCOUNT_EXPIRED (1793)
value ERROR_ACCOUNT_LOCKED_OUT (1909)
value ERROR_ACCOUNT_RESTRICTION (1327)
value ERROR_ACPI_ERROR (669)
value ERROR_ACTIVATION_COUNT_EXCEEDED (7059)
value ERROR_ACTIVE_CONNECTIONS (2402)
value ERROR_ADAP_HDW_ERR (57)
value ERROR_ADDRESS_ALREADY_ASSOCIATED (1227)
value ERROR_ADDRESS_NOT_ASSOCIATED (1228)
value ERROR_ADVANCED_INSTALLER_FAILED (14099)
value ERROR_ALERTED (739)
value ERROR_ALIAS_EXISTS (1379)
value ERROR_ALLOCATE_BUCKET (602)
value ERROR_ALLOTTED_SPACE_EXCEEDED (1344)
value ERROR_ALL_NODES_NOT_AVAILABLE (5037)
value ERROR_ALL_SIDS_FILTERED (_HRESULT_TYPEDEF_(0xC0090002L))
value ERROR_ALL_USER_TRUST_QUOTA_EXCEEDED (1933)
value ERROR_ALREADY_ASSIGNED (85)
value ERROR_ALREADY_EXISTS (183)
value ERROR_ALREADY_FIBER (1280)
value ERROR_ALREADY_HAS_STREAM_ID (4444)
value ERROR_ALREADY_INITIALIZED (1247)
value ERROR_ALREADY_REGISTERED (1242)
value ERROR_ALREADY_RUNNING_LKG (1074)
value ERROR_ALREADY_THREAD (1281)
value ERROR_ALREADY_WAITING (1904)
value ERROR_AMBIGUOUS_SYSTEM_DEVICE (15250)
value ERROR_API_UNAVAILABLE (15841)
value ERROR_APPCONTAINER_REQUIRED (4251)
value ERROR_APPEXEC_APP_COMPAT_BLOCK (3068)
value ERROR_APPEXEC_CALLER_WAIT_TIMEOUT (3069)
value ERROR_APPEXEC_CALLER_WAIT_TIMEOUT_LICENSING (3071)
value ERROR_APPEXEC_CALLER_WAIT_TIMEOUT_RESOURCES (3072)
value ERROR_APPEXEC_CALLER_WAIT_TIMEOUT_TERMINATION (3070)
value ERROR_APPEXEC_CONDITION_NOT_SATISFIED (3060)
value ERROR_APPEXEC_HANDLE_INVALIDATED (3061)
value ERROR_APPEXEC_HOST_ID_MISMATCH (3066)
value ERROR_APPEXEC_INVALID_HOST_GENERATION (3062)
value ERROR_APPEXEC_INVALID_HOST_STATE (3064)
value ERROR_APPEXEC_NO_DONOR (3065)
value ERROR_APPEXEC_UNEXPECTED_PROCESS_REGISTRATION (3063)
value ERROR_APPEXEC_UNKNOWN_USER (3067)
value ERROR_APPHELP_BLOCK (1259)
value ERROR_APPINSTALLER_ACTIVATION_BLOCKED (15646)
value ERROR_APPINSTALLER_IS_MANAGED_BY_SYSTEM (15672)
value ERROR_APPINSTALLER_URI_IN_USE (15671)
value ERROR_APPX_FILE_NOT_ENCRYPTED (409)
value ERROR_APPX_INTEGRITY_FAILURE_CLR_NGEN (15624)
value ERROR_APPX_RAW_DATA_WRITE_FAILED (15648)
value ERROR_APP_DATA_CORRUPT (4402)
value ERROR_APP_DATA_EXPIRED (4401)
value ERROR_APP_DATA_LIMIT_EXCEEDED (4403)
value ERROR_APP_DATA_NOT_FOUND (4400)
value ERROR_APP_DATA_REBOOT_REQUIRED (4404)
value ERROR_APP_HANG (1298)
value ERROR_APP_INIT_FAILURE (575)
value ERROR_APP_WRONG_OS (1151)
value ERROR_ARBITRATION_UNHANDLED (723)
value ERROR_ARENA_TRASHED (7)
value ERROR_ARITHMETIC_OVERFLOW (534)
value ERROR_ASSERTION_FAILURE (668)
value ERROR_ATOMIC_LOCKS_NOT_SUPPORTED (174)
value ERROR_ATTRIBUTE_NOT_PRESENT (_HRESULT_TYPEDEF_(0x8083000AL))
value ERROR_AUDITING_DISABLED (_HRESULT_TYPEDEF_(0xC0090001L))
value ERROR_AUDIT_FAILED (606)
value ERROR_AUTHENTICATION_FIREWALL_FAILED (1935)
value ERROR_AUTHIP_FAILURE (1469)
value ERROR_BACKUP_CONTROLLER (586)
value ERROR_BADDB (1009)
value ERROR_BADKEY (1010)
value ERROR_BADSTARTPOSITION (778)
value ERROR_BAD_ACCESSOR_FLAGS (773)
value ERROR_BAD_ARGUMENTS (160)
value ERROR_BAD_CLUSTERS (6849)
value ERROR_BAD_COMMAND (22)
value ERROR_BAD_COMPRESSION_BUFFER (605)
value ERROR_BAD_CONFIGURATION (1610)
value ERROR_BAD_CURRENT_DIRECTORY (703)
value ERROR_BAD_DESCRIPTOR_FORMAT (1361)
value ERROR_BAD_DEVICE (1200)
value ERROR_BAD_DEVICE_PATH (330)
value ERROR_BAD_DEV_TYPE (66)
value ERROR_BAD_DLL_ENTRYPOINT (609)
value ERROR_BAD_DRIVER (2001)
value ERROR_BAD_DRIVER_LEVEL (119)
value ERROR_BAD_ENVIRONMENT (10)
value ERROR_BAD_EXE_FORMAT (193)
value ERROR_BAD_FILE_TYPE (222)
value ERROR_BAD_FORMAT (11)
value ERROR_BAD_FUNCTION_TABLE (559)
value ERROR_BAD_IMPERSONATION_LEVEL (1346)
value ERROR_BAD_INHERITANCE_ACL (1340)
value ERROR_BAD_LENGTH (24)
value ERROR_BAD_LOGON_SESSION_STATE (1365)
value ERROR_BAD_MCFG_TABLE (791)
value ERROR_BAD_NETPATH (53)
value ERROR_BAD_NET_NAME (67)
value ERROR_BAD_NET_RESP (58)
value ERROR_BAD_PATHNAME (161)
value ERROR_BAD_PIPE (230)
value ERROR_BAD_PROFILE (1206)
value ERROR_BAD_PROVIDER (1204)
value ERROR_BAD_QUERY_SYNTAX (1615)
value ERROR_BAD_RECOVERY_POLICY (6012)
value ERROR_BAD_REM_ADAP (60)
value ERROR_BAD_SERVICE_ENTRYPOINT (610)
value ERROR_BAD_STACK (543)
value ERROR_BAD_THREADID_ADDR (159)
value ERROR_BAD_TOKEN_TYPE (1349)
value ERROR_BAD_UNIT (20)
value ERROR_BAD_USERNAME (2202)
value ERROR_BAD_USER_PROFILE (1253)
value ERROR_BAD_VALIDATION_CLASS (1348)
value ERROR_BCD_NOT_ALL_ENTRIES_IMPORTED (_NDIS_ERROR_TYPEDEF_(0x80390001L))
value ERROR_BCD_NOT_ALL_ENTRIES_SYNCHRONIZED (_NDIS_ERROR_TYPEDEF_(0x80390003L))
value ERROR_BCD_TOO_MANY_ELEMENTS (_NDIS_ERROR_TYPEDEF_(0xC0390002L))
value ERROR_BEGINNING_OF_MEDIA (1102)
value ERROR_BEYOND_VDL (1289)
value ERROR_BIDI_DEVICE_CONFIG_UNCHANGED ((ERROR_BIDI_ERROR_BASE + 14))
value ERROR_BIDI_DEVICE_OFFLINE ((ERROR_BIDI_ERROR_BASE + 4))
value ERROR_BIDI_ERROR_BASE (13000)
value ERROR_BIDI_GET_ARGUMENT_NOT_SUPPORTED ((ERROR_BIDI_ERROR_BASE + 12))
value ERROR_BIDI_GET_MISSING_ARGUMENT ((ERROR_BIDI_ERROR_BASE + 13))
value ERROR_BIDI_GET_REQUIRES_ARGUMENT ((ERROR_BIDI_ERROR_BASE + 11))
value ERROR_BIDI_NOT_SUPPORTED (ERROR_NOT_SUPPORTED)
value ERROR_BIDI_NO_BIDI_SCHEMA_EXTENSIONS ((ERROR_BIDI_ERROR_BASE + 16))
value ERROR_BIDI_NO_LOCALIZED_RESOURCES ((ERROR_BIDI_ERROR_BASE + 15))
value ERROR_BIDI_SCHEMA_NOT_SUPPORTED ((ERROR_BIDI_ERROR_BASE + 5))
value ERROR_BIDI_SCHEMA_READ_ONLY ((ERROR_BIDI_ERROR_BASE + 2))
value ERROR_BIDI_SCHEMA_WRITE_ONLY ((ERROR_BIDI_ERROR_BASE + 10))
value ERROR_BIDI_SERVER_OFFLINE ((ERROR_BIDI_ERROR_BASE + 3))
value ERROR_BIDI_SET_DIFFERENT_TYPE ((ERROR_BIDI_ERROR_BASE + 6))
value ERROR_BIDI_SET_INVALID_SCHEMAPATH ((ERROR_BIDI_ERROR_BASE + 8))
value ERROR_BIDI_SET_MULTIPLE_SCHEMAPATH ((ERROR_BIDI_ERROR_BASE + 7))
value ERROR_BIDI_SET_UNKNOWN_FAILURE ((ERROR_BIDI_ERROR_BASE + 9))
value ERROR_BIDI_STATUS_OK (0)
value ERROR_BIDI_STATUS_WARNING ((ERROR_BIDI_ERROR_BASE + 1))
value ERROR_BIDI_UNSUPPORTED_CLIENT_LANGUAGE ((ERROR_BIDI_ERROR_BASE + 17))
value ERROR_BIDI_UNSUPPORTED_RESOURCE_FORMAT ((ERROR_BIDI_ERROR_BASE + 18))
value ERROR_BIOS_FAILED_TO_CONNECT_INTERRUPT (585)
value ERROR_BIZRULES_NOT_ENABLED (_HRESULT_TYPEDEF_(0xC0090003L))
value ERROR_BLOCKED_BY_PARENTAL_CONTROLS (346)
value ERROR_BLOCK_SHARED (514)
value ERROR_BLOCK_SOURCE_WEAK_REFERENCE_INVALID (512)
value ERROR_BLOCK_TARGET_WEAK_REFERENCE_INVALID (513)
value ERROR_BLOCK_TOO_MANY_REFERENCES (347)
value ERROR_BLOCK_WEAK_REFERENCE_INVALID (511)
value ERROR_BOOT_ALREADY_ACCEPTED (1076)
value ERROR_BROKEN_PIPE (109)
value ERROR_BUFFER_ALL_ZEROS (754)
value ERROR_BUFFER_OVERFLOW (111)
value ERROR_BUSY (170)
value ERROR_BUSY_DRIVE (142)
value ERROR_BUS_RESET (1111)
value ERROR_BYPASSIO_FLT_NOT_SUPPORTED (506)
value ERROR_CACHE_PAGE_LOCKED (752)
value ERROR_CALLBACK_INVOKE_INLINE (812)
value ERROR_CALLBACK_POP_STACK (768)
value ERROR_CALLBACK_SUPPLIED_INVALID_DATA (1273)
value ERROR_CALL_NOT_IMPLEMENTED (120)
value ERROR_CANCELLED (1223)
value ERROR_CANCEL_VIOLATION (173)
value ERROR_CANNOT_ABORT_TRANSACTIONS (6848)
value ERROR_CANNOT_ACCEPT_TRANSACTED_WORK (6847)
value ERROR_CANNOT_BREAK_OPLOCK (802)
value ERROR_CANNOT_COPY (266)
value ERROR_CANNOT_DETECT_DRIVER_FAILURE (1080)
value ERROR_CANNOT_DETECT_PROCESS_ABORT (1081)
value ERROR_CANNOT_EXECUTE_FILE_IN_TRANSACTION (6838)
value ERROR_CANNOT_FIND_WND_CLASS (1407)
value ERROR_CANNOT_GRANT_REQUESTED_OPLOCK (801)
value ERROR_CANNOT_IMPERSONATE (1368)
value ERROR_CANNOT_LOAD_REGISTRY_FILE (589)
value ERROR_CANNOT_MAKE (82)
value ERROR_CANNOT_OPEN_PROFILE (1205)
value ERROR_CANNOT_SWITCH_RUNLEVEL (15400)
value ERROR_CANTFETCHBACKWARDS (770)
value ERROR_CANTOPEN (1011)
value ERROR_CANTREAD (1012)
value ERROR_CANTSCROLLBACKWARDS (771)
value ERROR_CANTWRITE (1013)
value ERROR_CANT_ACCESS_DOMAIN_INFO (1351)
value ERROR_CANT_ACCESS_FILE (1920)
value ERROR_CANT_BREAK_TRANSACTIONAL_DEPENDENCY (6824)
value ERROR_CANT_CLEAR_ENCRYPTION_FLAG (432)
value ERROR_CANT_CREATE_MORE_STREAM_MINIVERSIONS (6812)
value ERROR_CANT_CROSS_RM_BOUNDARY (6825)
value ERROR_CANT_DELETE_LAST_ITEM (4335)
value ERROR_CANT_DISABLE_MANDATORY (1310)
value ERROR_CANT_ENABLE_DENY_ONLY (629)
value ERROR_CANT_EVICT_ACTIVE_NODE (5009)
value ERROR_CANT_OPEN_ANONYMOUS (1347)
value ERROR_CANT_OPEN_MINIVERSION_WITH_MODIFY_INTENT (6811)
value ERROR_CANT_RECOVER_WITH_HANDLE_OPEN (6818)
value ERROR_CANT_RESOLVE_FILENAME (1921)
value ERROR_CANT_TERMINATE_SELF (555)
value ERROR_CANT_WAIT (554)
value ERROR_CAN_NOT_COMPLETE (1003)
value ERROR_CAN_NOT_DEL_LOCAL_WINS (4001)
value ERROR_CAPAUTHZ_CHANGE_TYPE (451)
value ERROR_CAPAUTHZ_DB_CORRUPTED (455)
value ERROR_CAPAUTHZ_NOT_AUTHORIZED (453)
value ERROR_CAPAUTHZ_NOT_DEVUNLOCKED (450)
value ERROR_CAPAUTHZ_NOT_PROVISIONED (452)
value ERROR_CAPAUTHZ_NO_POLICY (454)
value ERROR_CAPAUTHZ_SCCD_DEV_MODE_REQUIRED (459)
value ERROR_CAPAUTHZ_SCCD_INVALID_CATALOG (456)
value ERROR_CAPAUTHZ_SCCD_NO_AUTH_ENTITY (457)
value ERROR_CAPAUTHZ_SCCD_NO_CAPABILITY_MATCH (460)
value ERROR_CAPAUTHZ_SCCD_PARSE_ERROR (458)
value ERROR_CARDBUS_NOT_SUPPORTED (724)
value ERROR_CASE_DIFFERING_NAMES_IN_DIR (424)
value ERROR_CASE_SENSITIVE_PATH (442)
value ERROR_CERTIFICATE_VALIDATION_PREFERENCE_CONFLICT (817)
value ERROR_CHECKING_FILE_SYSTEM (712)
value ERROR_CHECKOUT_REQUIRED (221)
value ERROR_CHILD_MUST_BE_VOLATILE (1021)
value ERROR_CHILD_NOT_COMPLETE (129)
value ERROR_CHILD_PROCESS_BLOCKED (367)
value ERROR_CHILD_WINDOW_MENU (1436)
value ERROR_CIMFS_IMAGE_CORRUPT (470)
value ERROR_CIMFS_IMAGE_VERSION_NOT_SUPPORTED (471)
value ERROR_CIRCULAR_DEPENDENCY (1059)
value ERROR_CLASSIC_COMPAT_MODE_NOT_ALLOWED (15667)
value ERROR_CLASS_ALREADY_EXISTS (1410)
value ERROR_CLASS_DOES_NOT_EXIST (1411)
value ERROR_CLASS_HAS_WINDOWS (1412)
value ERROR_CLEANER_CARTRIDGE_INSTALLED (4340)
value ERROR_CLEANER_CARTRIDGE_SPENT (4333)
value ERROR_CLEANER_SLOT_NOT_SET (4332)
value ERROR_CLEANER_SLOT_SET (4331)
value ERROR_CLIENT_SERVER_PARAMETERS_INVALID (597)
value ERROR_CLIPBOARD_NOT_OPEN (1418)
value ERROR_CLIPPING_NOT_SUPPORTED (2005)
value ERROR_CLIP_DEVICE_LICENSE_MISSING (_HRESULT_TYPEDEF_(0xC0EA0003L))
value ERROR_CLIP_KEYHOLDER_LICENSE_MISSING_OR_INVALID (_HRESULT_TYPEDEF_(0xC0EA0005L))
value ERROR_CLIP_LICENSE_DEVICE_ID_MISMATCH (_HRESULT_TYPEDEF_(0xC0EA000AL))
value ERROR_CLIP_LICENSE_EXPIRED (_HRESULT_TYPEDEF_(0xC0EA0006L))
value ERROR_CLIP_LICENSE_HARDWARE_ID_OUT_OF_TOLERANCE (_HRESULT_TYPEDEF_(0xC0EA0009L))
value ERROR_CLIP_LICENSE_INVALID_SIGNATURE (_HRESULT_TYPEDEF_(0xC0EA0004L))
value ERROR_CLIP_LICENSE_NOT_FOUND (_HRESULT_TYPEDEF_(0xC0EA0002L))
value ERROR_CLIP_LICENSE_NOT_SIGNED (_HRESULT_TYPEDEF_(0xC0EA0008L))
value ERROR_CLIP_LICENSE_SIGNED_BY_UNKNOWN_SOURCE (_HRESULT_TYPEDEF_(0xC0EA0007L))
value ERROR_CLOUD_FILE_ACCESS_DENIED (395)
value ERROR_CLOUD_FILE_ALREADY_CONNECTED (378)
value ERROR_CLOUD_FILE_AUTHENTICATION_FAILED (386)
value ERROR_CLOUD_FILE_CONNECTED_PROVIDER_ONLY (382)
value ERROR_CLOUD_FILE_DEHYDRATION_DISALLOWED (434)
value ERROR_CLOUD_FILE_INCOMPATIBLE_HARDLINKS (396)
value ERROR_CLOUD_FILE_INSUFFICIENT_RESOURCES (387)
value ERROR_CLOUD_FILE_INVALID_REQUEST (380)
value ERROR_CLOUD_FILE_IN_USE (391)
value ERROR_CLOUD_FILE_METADATA_CORRUPT (363)
value ERROR_CLOUD_FILE_METADATA_TOO_LARGE (364)
value ERROR_CLOUD_FILE_NETWORK_UNAVAILABLE (388)
value ERROR_CLOUD_FILE_NOT_IN_SYNC (377)
value ERROR_CLOUD_FILE_NOT_SUPPORTED (379)
value ERROR_CLOUD_FILE_NOT_UNDER_SYNC_ROOT (390)
value ERROR_CLOUD_FILE_PINNED (392)
value ERROR_CLOUD_FILE_PROPERTY_BLOB_CHECKSUM_MISMATCH (366)
value ERROR_CLOUD_FILE_PROPERTY_BLOB_TOO_LARGE (365)
value ERROR_CLOUD_FILE_PROPERTY_CORRUPT (394)
value ERROR_CLOUD_FILE_PROPERTY_LOCK_CONFLICT (397)
value ERROR_CLOUD_FILE_PROPERTY_VERSION_NOT_SUPPORTED (375)
value ERROR_CLOUD_FILE_PROVIDER_NOT_RUNNING (362)
value ERROR_CLOUD_FILE_PROVIDER_TERMINATED (404)
value ERROR_CLOUD_FILE_READ_ONLY_VOLUME (381)
value ERROR_CLOUD_FILE_REQUEST_ABORTED (393)
value ERROR_CLOUD_FILE_REQUEST_CANCELED (398)
value ERROR_CLOUD_FILE_REQUEST_TIMEOUT (426)
value ERROR_CLOUD_FILE_SYNC_ROOT_METADATA_CORRUPT (358)
value ERROR_CLOUD_FILE_TOO_MANY_PROPERTY_BLOBS (374)
value ERROR_CLOUD_FILE_UNSUCCESSFUL (389)
value ERROR_CLOUD_FILE_US_MESSAGE_TIMEOUT (475)
value ERROR_CLOUD_FILE_VALIDATION_FAILED (383)
value ERROR_CLUSCFG_ALREADY_COMMITTED (5901)
value ERROR_CLUSCFG_ROLLBACK_FAILED (5902)
value ERROR_CLUSCFG_SYSTEM_DISK_DRIVE_LETTER_CONFLICT (5903)
value ERROR_CLUSTERLOG_CHKPOINT_NOT_FOUND (5032)
value ERROR_CLUSTERLOG_CORRUPT (5029)
value ERROR_CLUSTERLOG_EXCEEDS_MAXSIZE (5031)
value ERROR_CLUSTERLOG_NOT_ENOUGH_SPACE (5033)
value ERROR_CLUSTERLOG_RECORD_EXCEEDS_MAXSIZE (5030)
value ERROR_CLUSTERSET_MANAGEMENT_CLUSTER_UNREACHABLE (5999)
value ERROR_CLUSTER_AFFINITY_CONFLICT (5971)
value ERROR_CLUSTER_BACKUP_IN_PROGRESS (5949)
value ERROR_CLUSTER_CANNOT_RETURN_PROPERTIES (5968)
value ERROR_CLUSTER_CANT_CREATE_DUP_CLUSTER_NAME (5900)
value ERROR_CLUSTER_CANT_DESERIALIZE_DATA (5923)
value ERROR_CLUSTER_CSV_INVALID_HANDLE (5989)
value ERROR_CLUSTER_CSV_IO_PAUSE_TIMEOUT (5979)
value ERROR_CLUSTER_CSV_SUPPORTED_ONLY_ON_COORDINATOR (5990)
value ERROR_CLUSTER_DATABASE_SEQMISMATCH (5083)
value ERROR_CLUSTER_DATABASE_TRANSACTION_IN_PROGRESS (5918)
value ERROR_CLUSTER_DATABASE_TRANSACTION_NOT_IN_PROGRESS (5919)
value ERROR_CLUSTER_DATABASE_UPDATE_CONDITION_FAILED (5986)
value ERROR_CLUSTER_DISK_NOT_CONNECTED (5963)
value ERROR_CLUSTER_EVICT_INVALID_REQUEST (5939)
value ERROR_CLUSTER_EVICT_WITHOUT_CLEANUP (5896)
value ERROR_CLUSTER_FAULT_DOMAIN_INVALID_HIERARCHY (5995)
value ERROR_CLUSTER_FAULT_DOMAIN_PARENT_NOT_FOUND (5994)
value ERROR_CLUSTER_GROUP_BUSY (5944)
value ERROR_CLUSTER_GROUP_MOVING (5908)
value ERROR_CLUSTER_GROUP_QUEUED (5959)
value ERROR_CLUSTER_GROUP_SINGLETON_RESOURCE (5941)
value ERROR_CLUSTER_GUM_NOT_LOCKER (5085)
value ERROR_CLUSTER_INCOMPATIBLE_VERSIONS (5075)
value ERROR_CLUSTER_INSTANCE_ID_MISMATCH (5893)
value ERROR_CLUSTER_INTERNAL_INVALID_FUNCTION (5912)
value ERROR_CLUSTER_INVALID_INFRASTRUCTURE_FILESERVER_NAME (5998)
value ERROR_CLUSTER_INVALID_NETWORK (5054)
value ERROR_CLUSTER_INVALID_NETWORK_PROVIDER (5049)
value ERROR_CLUSTER_INVALID_NODE (5039)
value ERROR_CLUSTER_INVALID_NODE_WEIGHT (5954)
value ERROR_CLUSTER_INVALID_REQUEST (5048)
value ERROR_CLUSTER_INVALID_SECURITY_DESCRIPTOR (5946)
value ERROR_CLUSTER_INVALID_STRING_FORMAT (5917)
value ERROR_CLUSTER_INVALID_STRING_TERMINATION (5916)
value ERROR_CLUSTER_IPADDR_IN_USE (5057)
value ERROR_CLUSTER_JOIN_ABORTED (5074)
value ERROR_CLUSTER_JOIN_IN_PROGRESS (5041)
value ERROR_CLUSTER_JOIN_NOT_IN_PROGRESS (5053)
value ERROR_CLUSTER_LAST_INTERNAL_NETWORK (5066)
value ERROR_CLUSTER_LOCAL_NODE_NOT_FOUND (5043)
value ERROR_CLUSTER_MAXNUM_OF_RESOURCES_EXCEEDED (5076)
value ERROR_CLUSTER_MAX_NODES_IN_CLUSTER (5934)
value ERROR_CLUSTER_MEMBERSHIP_HALT (5892)
value ERROR_CLUSTER_MEMBERSHIP_INVALID_STATE (5890)
value ERROR_CLUSTER_MISMATCHED_COMPUTER_ACCT_NAME (5905)
value ERROR_CLUSTER_NETINTERFACE_EXISTS (5046)
value ERROR_CLUSTER_NETINTERFACE_NOT_FOUND (5047)
value ERROR_CLUSTER_NETWORK_ALREADY_OFFLINE (5064)
value ERROR_CLUSTER_NETWORK_ALREADY_ONLINE (5063)
value ERROR_CLUSTER_NETWORK_EXISTS (5044)
value ERROR_CLUSTER_NETWORK_HAS_DEPENDENTS (5067)
value ERROR_CLUSTER_NETWORK_NOT_FOUND (5045)
value ERROR_CLUSTER_NETWORK_NOT_FOUND_FOR_IP (5894)
value ERROR_CLUSTER_NETWORK_NOT_INTERNAL (5060)
value ERROR_CLUSTER_NODE_ALREADY_DOWN (5062)
value ERROR_CLUSTER_NODE_ALREADY_HAS_DFS_ROOT (5088)
value ERROR_CLUSTER_NODE_ALREADY_MEMBER (5065)
value ERROR_CLUSTER_NODE_ALREADY_UP (5061)
value ERROR_CLUSTER_NODE_DOWN (5050)
value ERROR_CLUSTER_NODE_DRAIN_IN_PROGRESS (5962)
value ERROR_CLUSTER_NODE_EXISTS (5040)
value ERROR_CLUSTER_NODE_IN_GRACE_PERIOD (5978)
value ERROR_CLUSTER_NODE_ISOLATED (5984)
value ERROR_CLUSTER_NODE_NOT_FOUND (5042)
value ERROR_CLUSTER_NODE_NOT_MEMBER (5052)
value ERROR_CLUSTER_NODE_NOT_PAUSED (5058)
value ERROR_CLUSTER_NODE_NOT_READY (5072)
value ERROR_CLUSTER_NODE_PAUSED (5070)
value ERROR_CLUSTER_NODE_QUARANTINED (5985)
value ERROR_CLUSTER_NODE_SHUTTING_DOWN (5073)
value ERROR_CLUSTER_NODE_UNREACHABLE (5051)
value ERROR_CLUSTER_NODE_UP (5056)
value ERROR_CLUSTER_NOT_INSTALLED (5932)
value ERROR_CLUSTER_NOT_SHARED_VOLUME (5945)
value ERROR_CLUSTER_NO_NET_ADAPTERS (5906)
value ERROR_CLUSTER_NO_QUORUM (5925)
value ERROR_CLUSTER_NO_RPC_PACKAGES_REGISTERED (5081)
value ERROR_CLUSTER_NO_SECURITY_CONTEXT (5059)
value ERROR_CLUSTER_NULL_DATA (5920)
value ERROR_CLUSTER_OBJECT_ALREADY_USED (5936)
value ERROR_CLUSTER_OBJECT_IS_CLUSTER_SET_VM (6250)
value ERROR_CLUSTER_OLD_VERSION (5904)
value ERROR_CLUSTER_OWNER_NOT_IN_PREFLIST (5082)
value ERROR_CLUSTER_PARAMETER_MISMATCH (5897)
value ERROR_CLUSTER_PARAMETER_OUT_OF_BOUNDS (5913)
value ERROR_CLUSTER_PARTIAL_READ (5921)
value ERROR_CLUSTER_PARTIAL_SEND (5914)
value ERROR_CLUSTER_PARTIAL_WRITE (5922)
value ERROR_CLUSTER_POISONED (5907)
value ERROR_CLUSTER_PROPERTY_DATA_TYPE_MISMATCH (5895)
value ERROR_CLUSTER_QUORUMLOG_NOT_FOUND (5891)
value ERROR_CLUSTER_REGISTRY_INVALID_FUNCTION (5915)
value ERROR_CLUSTER_RESNAME_NOT_FOUND (5080)
value ERROR_CLUSTER_RESOURCES_MUST_BE_ONLINE_ON_THE_SAME_NODE (5933)
value ERROR_CLUSTER_RESOURCE_CONFIGURATION_ERROR (5943)
value ERROR_CLUSTER_RESOURCE_CONTAINS_UNSUPPORTED_DIFF_AREA_FOR_SHARED_VOLUMES (5969)
value ERROR_CLUSTER_RESOURCE_DOES_NOT_SUPPORT_UNMONITORED (5982)
value ERROR_CLUSTER_RESOURCE_IS_IN_MAINTENANCE_MODE (5970)
value ERROR_CLUSTER_RESOURCE_IS_REPLICATED (5983)
value ERROR_CLUSTER_RESOURCE_IS_REPLICA_VIRTUAL_MACHINE (5972)
value ERROR_CLUSTER_RESOURCE_LOCKED_STATUS (5960)
value ERROR_CLUSTER_RESOURCE_NOT_MONITORED (5981)
value ERROR_CLUSTER_RESOURCE_PROVIDER_FAILED (5942)
value ERROR_CLUSTER_RESOURCE_TYPE_BUSY (5909)
value ERROR_CLUSTER_RESOURCE_TYPE_NOT_FOUND (5078)
value ERROR_CLUSTER_RESOURCE_VETOED_CALL (5955)
value ERROR_CLUSTER_RESOURCE_VETOED_MOVE_INCOMPATIBLE_NODES (5953)
value ERROR_CLUSTER_RESOURCE_VETOED_MOVE_NOT_ENOUGH_RESOURCES_ON_DESTINATION (5957)
value ERROR_CLUSTER_RESOURCE_VETOED_MOVE_NOT_ENOUGH_RESOURCES_ON_SOURCE (5958)
value ERROR_CLUSTER_RESTYPE_NOT_SUPPORTED (5079)
value ERROR_CLUSTER_RHS_FAILED_INITIALIZATION (5931)
value ERROR_CLUSTER_SHARED_VOLUMES_IN_USE (5947)
value ERROR_CLUSTER_SHARED_VOLUME_FAILOVER_NOT_ALLOWED (5961)
value ERROR_CLUSTER_SHARED_VOLUME_NOT_REDIRECTED (5967)
value ERROR_CLUSTER_SHARED_VOLUME_REDIRECTED (5966)
value ERROR_CLUSTER_SHUTTING_DOWN (5022)
value ERROR_CLUSTER_SINGLETON_RESOURCE (5940)
value ERROR_CLUSTER_SPACE_DEGRADED (5987)
value ERROR_CLUSTER_SYSTEM_CONFIG_CHANGED (5077)
value ERROR_CLUSTER_TOKEN_DELEGATION_NOT_SUPPORTED (5988)
value ERROR_CLUSTER_TOO_MANY_NODES (5935)
value ERROR_CLUSTER_UPGRADE_FIX_QUORUM_NOT_SUPPORTED (5974)
value ERROR_CLUSTER_UPGRADE_INCOMPATIBLE_VERSIONS (5973)
value ERROR_CLUSTER_UPGRADE_INCOMPLETE (5977)
value ERROR_CLUSTER_UPGRADE_IN_PROGRESS (5976)
value ERROR_CLUSTER_UPGRADE_RESTART_REQUIRED (5975)
value ERROR_CLUSTER_USE_SHARED_VOLUMES_API (5948)
value ERROR_CLUSTER_WATCHDOG_TERMINATING (5952)
value ERROR_CLUSTER_WRONG_OS_VERSION (5899)
value ERROR_COLORSPACE_MISMATCH (2021)
value ERROR_COMMITMENT_LIMIT (1455)
value ERROR_COMMITMENT_MINIMUM (635)
value ERROR_COMPRESSED_FILE_NOT_SUPPORTED (335)
value ERROR_COMPRESSION_DISABLED (769)
value ERROR_COMPRESSION_NOT_ALLOWED_IN_TRANSACTION (6850)
value ERROR_COMPRESSION_NOT_BENEFICIAL (344)
value ERROR_COM_TASK_STOP_PENDING (15501)
value ERROR_CONNECTED_OTHER_PASSWORD (2108)
value ERROR_CONNECTED_OTHER_PASSWORD_DEFAULT (2109)
value ERROR_CONNECTION_ABORTED (1236)
value ERROR_CONNECTION_ACTIVE (1230)
value ERROR_CONNECTION_COUNT_LIMIT (1238)
value ERROR_CONNECTION_INVALID (1229)
value ERROR_CONNECTION_REFUSED (1225)
value ERROR_CONNECTION_UNAVAIL (1201)
value ERROR_CONTAINER_ASSIGNED (1504)
value ERROR_CONTENT_BLOCKED (1296)
value ERROR_CONTEXT_EXPIRED (1931)
value ERROR_CONTINUE (1246)
value ERROR_CONTROLLING_IEPORT (4329)
value ERROR_CONTROL_C_EXIT (572)
value ERROR_CONTROL_ID_NOT_FOUND (1421)
value ERROR_CONVERT_TO_LARGE (600)
value ERROR_CORE_DRIVER_PACKAGE_NOT_FOUND (3016)
value ERROR_CORE_RESOURCE (5026)
value ERROR_CORRUPT_LOG_CLEARED (798)
value ERROR_CORRUPT_LOG_CORRUPTED (795)
value ERROR_CORRUPT_LOG_DELETED_FULL (797)
value ERROR_CORRUPT_LOG_OVERFULL (794)
value ERROR_CORRUPT_LOG_UNAVAILABLE (796)
value ERROR_CORRUPT_SYSTEM_FILE (634)
value ERROR_COULD_NOT_INTERPRET (552)
value ERROR_COULD_NOT_RESIZE_LOG (6629)
value ERROR_COUNTER_TIMEOUT (1121)
value ERROR_CPU_SET_INVALID (813)
value ERROR_CRASH_DUMP (753)
value ERROR_CRC (23)
value ERROR_CREATE_FAILED (1631)
value ERROR_CRED_REQUIRES_CONFIRMATION (_HRESULT_TYPEDEF_(0x80097019L))
value ERROR_CRM_PROTOCOL_ALREADY_EXISTS (6710)
value ERROR_CRM_PROTOCOL_NOT_FOUND (6712)
value ERROR_CROSS_PARTITION_VIOLATION (1661)
value ERROR_CSCSHARE_OFFLINE (1262)
value ERROR_CSV_VOLUME_NOT_LOCAL (5951)
value ERROR_CS_ENCRYPTION_EXISTING_ENCRYPTED_FILE (6019)
value ERROR_CS_ENCRYPTION_FILE_NOT_CSE (6021)
value ERROR_CS_ENCRYPTION_INVALID_SERVER_RESPONSE (6017)
value ERROR_CS_ENCRYPTION_NEW_ENCRYPTED_FILE (6020)
value ERROR_CS_ENCRYPTION_UNSUPPORTED_SERVER (6018)
value ERROR_CTLOG_INCONSISTENT_TRACKING_FILE (_NDIS_ERROR_TYPEDEF_(0xC03A0024L))
value ERROR_CTLOG_INVALID_TRACKING_STATE (_NDIS_ERROR_TYPEDEF_(0xC03A0023L))
value ERROR_CTLOG_LOGFILE_SIZE_EXCEEDED_MAXSIZE (_NDIS_ERROR_TYPEDEF_(0xC03A0021L))
value ERROR_CTLOG_TRACKING_NOT_INITIALIZED (_NDIS_ERROR_TYPEDEF_(0xC03A0020L))
value ERROR_CTLOG_VHD_CHANGED_OFFLINE (_NDIS_ERROR_TYPEDEF_(0xC03A0022L))
value ERROR_CTX_ACCOUNT_RESTRICTION (7064)
value ERROR_CTX_BAD_VIDEO_MODE (7025)
value ERROR_CTX_CANNOT_MAKE_EVENTLOG_ENTRY (7005)
value ERROR_CTX_CDM_CONNECT (7066)
value ERROR_CTX_CDM_DISCONNECT (7067)
value ERROR_CTX_CLIENT_LICENSE_IN_USE (7052)
value ERROR_CTX_CLIENT_LICENSE_NOT_SET (7053)
value ERROR_CTX_CLIENT_QUERY_TIMEOUT (7040)
value ERROR_CTX_CLOSE_PENDING (7007)
value ERROR_CTX_CONSOLE_CONNECT (7042)
value ERROR_CTX_CONSOLE_DISCONNECT (7041)
value ERROR_CTX_ENCRYPTION_LEVEL_REQUIRED (7061)
value ERROR_CTX_GRAPHICS_INVALID (7035)
value ERROR_CTX_INVALID_MODEMNAME (7010)
value ERROR_CTX_INVALID_PD (7002)
value ERROR_CTX_INVALID_WD (7049)
value ERROR_CTX_LICENSE_CLIENT_INVALID (7055)
value ERROR_CTX_LICENSE_EXPIRED (7056)
value ERROR_CTX_LICENSE_NOT_AVAILABLE (7054)
value ERROR_CTX_LOGON_DISABLED (7037)
value ERROR_CTX_MODEM_INF_NOT_FOUND (7009)
value ERROR_CTX_MODEM_RESPONSE_BUSY (7015)
value ERROR_CTX_MODEM_RESPONSE_ERROR (7011)
value ERROR_CTX_MODEM_RESPONSE_NO_CARRIER (7013)
value ERROR_CTX_MODEM_RESPONSE_NO_DIALTONE (7014)
value ERROR_CTX_MODEM_RESPONSE_TIMEOUT (7012)
value ERROR_CTX_MODEM_RESPONSE_VOICE (7016)
value ERROR_CTX_NOT_CONSOLE (7038)
value ERROR_CTX_NO_FORCE_LOGOFF (7063)
value ERROR_CTX_NO_OUTBUF (7008)
value ERROR_CTX_PD_NOT_FOUND (7003)
value ERROR_CTX_SECURITY_LAYER_ERROR (7068)
value ERROR_CTX_SERVICE_NAME_COLLISION (7006)
value ERROR_CTX_SESSION_IN_USE (7062)
value ERROR_CTX_SHADOW_DENIED (7044)
value ERROR_CTX_SHADOW_DISABLED (7051)
value ERROR_CTX_SHADOW_ENDED_BY_MODE_CHANGE (7058)
value ERROR_CTX_SHADOW_INVALID (7050)
value ERROR_CTX_SHADOW_NOT_RUNNING (7057)
value ERROR_CTX_TD_ERROR (7017)
value ERROR_CTX_WD_NOT_FOUND (7004)
value ERROR_CTX_WINSTATIONS_DISABLED (7060)
value ERROR_CTX_WINSTATION_ACCESS_DENIED (7045)
value ERROR_CTX_WINSTATION_ALREADY_EXISTS (7023)
value ERROR_CTX_WINSTATION_BUSY (7024)
value ERROR_CTX_WINSTATION_NAME_INVALID (7001)
value ERROR_CTX_WINSTATION_NOT_FOUND (7022)
value ERROR_CURRENT_DIRECTORY (16)
value ERROR_CURRENT_DOMAIN_NOT_ALLOWED (1399)
value ERROR_CURRENT_TRANSACTION_NOT_VALID (6714)
value ERROR_DATABASE_BACKUP_CORRUPT (5087)
value ERROR_DATABASE_DOES_NOT_EXIST (1065)
value ERROR_DATABASE_FAILURE (4313)
value ERROR_DATABASE_FULL (4314)
value ERROR_DATATYPE_MISMATCH (1629)
value ERROR_DATA_CHECKSUM_ERROR (323)
value ERROR_DATA_LOST_REPAIR (6843)
value ERROR_DATA_NOT_ACCEPTED (592)
value ERROR_DAX_MAPPING_EXISTS (361)
value ERROR_DBG_ATTACH_PROCESS_FAILURE_LOCKDOWN (_HRESULT_TYPEDEF_(0x80B00002L))
value ERROR_DBG_COMMAND_EXCEPTION (697)
value ERROR_DBG_CONNECT_SERVER_FAILURE_LOCKDOWN (_HRESULT_TYPEDEF_(0x80B00003L))
value ERROR_DBG_CONTINUE (767)
value ERROR_DBG_CONTROL_BREAK (696)
value ERROR_DBG_CONTROL_C (693)
value ERROR_DBG_CREATE_PROCESS_FAILURE_LOCKDOWN (_HRESULT_TYPEDEF_(0x80B00001L))
value ERROR_DBG_EXCEPTION_HANDLED (766)
value ERROR_DBG_EXCEPTION_NOT_HANDLED (688)
value ERROR_DBG_PRINTEXCEPTION_C (694)
value ERROR_DBG_REPLY_LATER (689)
value ERROR_DBG_RIPEXCEPTION (695)
value ERROR_DBG_START_SERVER_FAILURE_LOCKDOWN (_HRESULT_TYPEDEF_(0x80B00004L))
value ERROR_DBG_TERMINATE_PROCESS (692)
value ERROR_DBG_TERMINATE_THREAD (691)
value ERROR_DBG_UNABLE_TO_PROVIDE_HANDLE (690)
value ERROR_DC_NOT_FOUND (1425)
value ERROR_DDE_FAIL (1156)
value ERROR_DEBUGGER_INACTIVE (1284)
value ERROR_DEBUG_ATTACH_FAILED (590)
value ERROR_DECRYPTION_FAILED (6001)
value ERROR_DELAY_LOAD_FAILED (1285)
value ERROR_DELETE_PENDING (303)
value ERROR_DELETING_EXISTING_APPLICATIONDATA_STORE_FAILED (15621)
value ERROR_DELETING_ICM_XFORM (2019)
value ERROR_DEPENDENCY_ALREADY_EXISTS (5003)
value ERROR_DEPENDENCY_NOT_ALLOWED (5069)
value ERROR_DEPENDENCY_NOT_FOUND (5002)
value ERROR_DEPENDENCY_TREE_TOO_COMPLEX (5929)
value ERROR_DEPENDENT_RESOURCE_EXISTS (5001)
value ERROR_DEPENDENT_RESOURCE_PROPERTY_CONFLICT (5924)
value ERROR_DEPENDENT_SERVICES_RUNNING (1051)
value ERROR_DEPLOYMENT_BLOCKED_BY_POLICY (15617)
value ERROR_DEPLOYMENT_BLOCKED_BY_PROFILE_POLICY (15651)
value ERROR_DEPLOYMENT_BLOCKED_BY_USER_LOG_OFF (15641)
value ERROR_DEPLOYMENT_BLOCKED_BY_VOLUME_POLICY_MACHINE (15650)
value ERROR_DEPLOYMENT_BLOCKED_BY_VOLUME_POLICY_PACKAGE (15649)
value ERROR_DEPLOYMENT_FAILED_CONFLICTING_MUTABLE_PACKAGE_DIRECTORY (15652)
value ERROR_DEPLOYMENT_OPTION_NOT_SUPPORTED (15645)
value ERROR_DESTINATION_ELEMENT_FULL (1161)
value ERROR_DESTROY_OBJECT_OF_OTHER_THREAD (1435)
value ERROR_DEVICE_ALREADY_ATTACHED (548)
value ERROR_DEVICE_ALREADY_REMEMBERED (1202)
value ERROR_DEVICE_DOOR_OPEN (1166)
value ERROR_DEVICE_ENUMERATION_ERROR (648)
value ERROR_DEVICE_FEATURE_NOT_SUPPORTED (316)
value ERROR_DEVICE_HARDWARE_ERROR (483)
value ERROR_DEVICE_HINT_NAME_BUFFER_TOO_SMALL (355)
value ERROR_DEVICE_IN_MAINTENANCE (359)
value ERROR_DEVICE_IN_USE (2404)
value ERROR_DEVICE_NOT_AVAILABLE (4319)
value ERROR_DEVICE_NOT_CONNECTED (1167)
value ERROR_DEVICE_NOT_PARTITIONED (1107)
value ERROR_DEVICE_NO_RESOURCES (322)
value ERROR_DEVICE_REINITIALIZATION_NEEDED (1164)
value ERROR_DEVICE_REMOVED (1617)
value ERROR_DEVICE_REQUIRES_CLEANING (1165)
value ERROR_DEVICE_RESET_REQUIRED (507)
value ERROR_DEVICE_SUPPORT_IN_PROGRESS (171)
value ERROR_DEVICE_UNREACHABLE (321)
value ERROR_DEV_NOT_EXIST (55)
value ERROR_DEV_SIDELOAD_LIMIT_EXCEEDED (15633)
value ERROR_DHCP_ADDRESS_CONFLICT (4100)
value ERROR_DIFFERENT_PROFILE_RESOURCE_MANAGER_EXIST (15144)
value ERROR_DIFFERENT_SERVICE_ACCOUNT (1079)
value ERROR_DIFFERENT_VERSION_OF_PACKAGED_SERVICE_INSTALLED (15654)
value ERROR_DIF_BINDING_API_NOT_FOUND (3199)
value ERROR_DIF_IOCALLBACK_NOT_REPLACED (3190)
value ERROR_DIF_LIVEDUMP_LIMIT_EXCEEDED (3191)
value ERROR_DIF_VOLATILE_DRIVER_HOTPATCHED (3193)
value ERROR_DIF_VOLATILE_DRIVER_IS_NOT_RUNNING (3195)
value ERROR_DIF_VOLATILE_INVALID_INFO (3194)
value ERROR_DIF_VOLATILE_NOT_ALLOWED (3198)
value ERROR_DIF_VOLATILE_PLUGIN_CHANGE_NOT_ALLOWED (3197)
value ERROR_DIF_VOLATILE_PLUGIN_IS_NOT_RUNNING (3196)
value ERROR_DIF_VOLATILE_SECTION_NOT_LOCKED (3192)
value ERROR_DIRECTORY (267)
value ERROR_DIRECTORY_NOT_RM (6803)
value ERROR_DIRECTORY_NOT_SUPPORTED (336)
value ERROR_DIRECT_ACCESS_HANDLE (130)
value ERROR_DIR_EFS_DISALLOWED (6010)
value ERROR_DIR_NOT_EMPTY (145)
value ERROR_DIR_NOT_ROOT (144)
value ERROR_DISCARDED (157)
value ERROR_DISK_CHANGE (107)
value ERROR_DISK_CORRUPT (1393)
value ERROR_DISK_FULL (112)
value ERROR_DISK_NOT_CSV_CAPABLE (5964)
value ERROR_DISK_OPERATION_FAILED (1127)
value ERROR_DISK_QUOTA_EXCEEDED (1295)
value ERROR_DISK_RECALIBRATE_FAILED (1126)
value ERROR_DISK_REPAIR_DISABLED (780)
value ERROR_DISK_REPAIR_REDIRECTED (792)
value ERROR_DISK_REPAIR_UNSUCCESSFUL (793)
value ERROR_DISK_RESET_FAILED (1128)
value ERROR_DISK_RESOURCES_EXHAUSTED (314)
value ERROR_DISK_TOO_FRAGMENTED (302)
value ERROR_DLL_INIT_FAILED (1114)
value ERROR_DLL_INIT_FAILED_LOGOFF (624)
value ERROR_DLL_MIGHT_BE_INCOMPATIBLE (687)
value ERROR_DLL_MIGHT_BE_INSECURE (686)
value ERROR_DLL_NOT_FOUND (1157)
value ERROR_DLP_POLICY_DENIES_OPERATION (446)
value ERROR_DLP_POLICY_SILENTLY_FAIL (449)
value ERROR_DLP_POLICY_WARNS_AGAINST_OPERATION (445)
value ERROR_DM_OPERATION_LIMIT_EXCEEDED (_HRESULT_TYPEDEF_(0xC0370600L))
value ERROR_DOMAIN_CONTROLLER_EXISTS (1250)
value ERROR_DOMAIN_CONTROLLER_NOT_FOUND (1908)
value ERROR_DOMAIN_CTRLR_CONFIG_ERROR (581)
value ERROR_DOMAIN_EXISTS (1356)
value ERROR_DOMAIN_LIMIT_EXCEEDED (1357)
value ERROR_DOMAIN_SID_SAME_AS_LOCAL_WORKSTATION (8644)
value ERROR_DOMAIN_TRUST_INCONSISTENT (1810)
value ERROR_DOWNGRADE_DETECTED (1265)
value ERROR_DPL_NOT_SUPPORTED_FOR_USER (423)
value ERROR_DRIVERS_LEAKING_LOCKED_PAGES (729)
value ERROR_DRIVER_BLOCKED (1275)
value ERROR_DRIVER_CANCEL_TIMEOUT (594)
value ERROR_DRIVER_DATABASE_ERROR (652)
value ERROR_DRIVER_FAILED_PRIOR_UNLOAD (654)
value ERROR_DRIVER_FAILED_SLEEP (633)
value ERROR_DRIVER_PROCESS_TERMINATED (1291)
value ERROR_DRIVE_LOCKED (108)
value ERROR_DRIVE_MEDIA_MISMATCH (4303)
value ERROR_DRIVE_NOT_INSTALLED (0x00000008)
value ERROR_DS_ADD_REPLICA_INHIBITED (8302)
value ERROR_DS_ADMIN_LIMIT_EXCEEDED (8228)
value ERROR_DS_AFFECTS_MULTIPLE_DSAS (8249)
value ERROR_DS_AG_CANT_HAVE_UNIVERSAL_MEMBER (8578)
value ERROR_DS_ALIASED_OBJ_MISSING (8334)
value ERROR_DS_ALIAS_DEREF_PROBLEM (8244)
value ERROR_DS_ALIAS_POINTS_TO_ALIAS (8336)
value ERROR_DS_ALIAS_PROBLEM (8241)
value ERROR_DS_ATTRIBUTE_OR_VALUE_EXISTS (8205)
value ERROR_DS_ATTRIBUTE_OWNED_BY_SAM (8346)
value ERROR_DS_ATTRIBUTE_TYPE_UNDEFINED (8204)
value ERROR_DS_ATT_ALREADY_EXISTS (8318)
value ERROR_DS_ATT_IS_NOT_ON_OBJ (8310)
value ERROR_DS_ATT_NOT_DEF_FOR_CLASS (8317)
value ERROR_DS_ATT_NOT_DEF_IN_SCHEMA (8303)
value ERROR_DS_ATT_SCHEMA_REQ_ID (8399)
value ERROR_DS_ATT_SCHEMA_REQ_SYNTAX (8416)
value ERROR_DS_ATT_VAL_ALREADY_EXISTS (8323)
value ERROR_DS_AUDIT_FAILURE (8625)
value ERROR_DS_AUTHORIZATION_FAILED (8599)
value ERROR_DS_AUTH_METHOD_NOT_SUPPORTED (8231)
value ERROR_DS_AUTH_UNKNOWN (8234)
value ERROR_DS_AUX_CLS_TEST_FAIL (8389)
value ERROR_DS_BACKLINK_WITHOUT_LINK (8482)
value ERROR_DS_BAD_ATT_SCHEMA_SYNTAX (8400)
value ERROR_DS_BAD_HIERARCHY_FILE (8425)
value ERROR_DS_BAD_INSTANCE_TYPE (8313)
value ERROR_DS_BAD_NAME_SYNTAX (8335)
value ERROR_DS_BAD_RDN_ATT_ID_SYNTAX (8392)
value ERROR_DS_BUILD_HIERARCHY_TABLE_FAILED (8426)
value ERROR_DS_BUSY (8206)
value ERROR_DS_CANT_ACCESS_REMOTE_PART_OF_AD (8585)
value ERROR_DS_CANT_ADD_ATT_VALUES (8320)
value ERROR_DS_CANT_ADD_SYSTEM_ONLY (8358)
value ERROR_DS_CANT_ADD_TO_GC (8550)
value ERROR_DS_CANT_CACHE_ATT (8401)
value ERROR_DS_CANT_CACHE_CLASS (8402)
value ERROR_DS_CANT_CREATE_IN_NONDOMAIN_NC (8553)
value ERROR_DS_CANT_CREATE_UNDER_SCHEMA (8510)
value ERROR_DS_CANT_DELETE (8398)
value ERROR_DS_CANT_DELETE_DSA_OBJ (8340)
value ERROR_DS_CANT_DEL_MASTER_CROSSREF (8375)
value ERROR_DS_CANT_DEMOTE_WITH_WRITEABLE_NC (8604)
value ERROR_DS_CANT_DEREF_ALIAS (8337)
value ERROR_DS_CANT_DERIVE_SPN_FOR_DELETED_DOMAIN (8603)
value ERROR_DS_CANT_DERIVE_SPN_WITHOUT_SERVER_REF (8589)
value ERROR_DS_CANT_FIND_DC_FOR_SRC_DOMAIN (8537)
value ERROR_DS_CANT_FIND_DSA_OBJ (8419)
value ERROR_DS_CANT_FIND_EXPECTED_NC (8420)
value ERROR_DS_CANT_FIND_NC_IN_CACHE (8421)
value ERROR_DS_CANT_MIX_MASTER_AND_REPS (8331)
value ERROR_DS_CANT_MOD_OBJ_CLASS (8215)
value ERROR_DS_CANT_MOD_PRIMARYGROUPID (8506)
value ERROR_DS_CANT_MOD_SYSTEM_ONLY (8369)
value ERROR_DS_CANT_MOVE_ACCOUNT_GROUP (8498)
value ERROR_DS_CANT_MOVE_APP_BASIC_GROUP (8608)
value ERROR_DS_CANT_MOVE_APP_QUERY_GROUP (8609)
value ERROR_DS_CANT_MOVE_DELETED_OBJECT (8489)
value ERROR_DS_CANT_MOVE_RESOURCE_GROUP (8499)
value ERROR_DS_CANT_ON_NON_LEAF (8213)
value ERROR_DS_CANT_ON_RDN (8214)
value ERROR_DS_CANT_REMOVE_ATT_CACHE (8403)
value ERROR_DS_CANT_REMOVE_CLASS_CACHE (8404)
value ERROR_DS_CANT_REM_MISSING_ATT (8324)
value ERROR_DS_CANT_REM_MISSING_ATT_VAL (8325)
value ERROR_DS_CANT_REPLACE_HIDDEN_REC (8424)
value ERROR_DS_CANT_RETRIEVE_ATTS (8481)
value ERROR_DS_CANT_RETRIEVE_CHILD (8422)
value ERROR_DS_CANT_RETRIEVE_DN (8405)
value ERROR_DS_CANT_RETRIEVE_INSTANCE (8407)
value ERROR_DS_CANT_RETRIEVE_SD (8526)
value ERROR_DS_CANT_START (8531)
value ERROR_DS_CANT_TREE_DELETE_CRITICAL_OBJ (8560)
value ERROR_DS_CANT_WITH_ACCT_GROUP_MEMBERSHPS (8493)
value ERROR_DS_CHILDREN_EXIST (8332)
value ERROR_DS_CLASS_MUST_BE_CONCRETE (8359)
value ERROR_DS_CLASS_NOT_DSA (8343)
value ERROR_DS_CLIENT_LOOP (8259)
value ERROR_DS_CODE_INCONSISTENCY (8408)
value ERROR_DS_COMPARE_FALSE (8229)
value ERROR_DS_COMPARE_TRUE (8230)
value ERROR_DS_CONFIDENTIALITY_REQUIRED (8237)
value ERROR_DS_CONFIG_PARAM_MISSING (8427)
value ERROR_DS_CONSTRAINT_VIOLATION (8239)
value ERROR_DS_CONSTRUCTED_ATT_MOD (8475)
value ERROR_DS_CONTROL_NOT_FOUND (8258)
value ERROR_DS_COULDNT_CONTACT_FSMO (8367)
value ERROR_DS_COULDNT_IDENTIFY_OBJECTS_FOR_TREE_DELETE (8503)
value ERROR_DS_COULDNT_LOCK_TREE_FOR_DELETE (8502)
value ERROR_DS_COULDNT_UPDATE_SPNS (8525)
value ERROR_DS_COUNTING_AB_INDICES_FAILED (8428)
value ERROR_DS_CROSS_DOMAIN_CLEANUP_REQD (8491)
value ERROR_DS_CROSS_DOM_MOVE_ERROR (8216)
value ERROR_DS_CROSS_NC_DN_RENAME (8368)
value ERROR_DS_CROSS_REF_BUSY (8602)
value ERROR_DS_CROSS_REF_EXISTS (8374)
value ERROR_DS_CR_IMPOSSIBLE_TO_VALIDATE (8495)
value ERROR_DS_DATABASE_ERROR (8409)
value ERROR_DS_DECODING_ERROR (8253)
value ERROR_DS_DESTINATION_AUDITING_NOT_ENABLED (8536)
value ERROR_DS_DESTINATION_DOMAIN_NOT_IN_FOREST (8535)
value ERROR_DS_DIFFERENT_REPL_EPOCHS (8593)
value ERROR_DS_DISALLOWED_IN_SYSTEM_CONTAINER (8615)
value ERROR_DS_DISALLOWED_NC_REDIRECT (8640)
value ERROR_DS_DNS_LOOKUP_FAILURE (8524)
value ERROR_DS_DOMAIN_NAME_EXISTS_IN_FOREST (8634)
value ERROR_DS_DOMAIN_RENAME_IN_PROGRESS (8612)
value ERROR_DS_DOMAIN_VERSION_TOO_HIGH (8564)
value ERROR_DS_DOMAIN_VERSION_TOO_LOW (8566)
value ERROR_DS_DRA_ABANDON_SYNC (8462)
value ERROR_DS_DRA_ACCESS_DENIED (8453)
value ERROR_DS_DRA_BAD_DN (8439)
value ERROR_DS_DRA_BAD_INSTANCE_TYPE (8445)
value ERROR_DS_DRA_BAD_NC (8440)
value ERROR_DS_DRA_BUSY (8438)
value ERROR_DS_DRA_CONNECTION_FAILED (8444)
value ERROR_DS_DRA_CORRUPT_UTD_VECTOR (8629)
value ERROR_DS_DRA_DB_ERROR (8451)
value ERROR_DS_DRA_DN_EXISTS (8441)
value ERROR_DS_DRA_EARLIER_SCHEMA_CONFLICT (8544)
value ERROR_DS_DRA_EXTN_CONNECTION_FAILED (8466)
value ERROR_DS_DRA_GENERIC (8436)
value ERROR_DS_DRA_INCOMPATIBLE_PARTIAL_SET (8464)
value ERROR_DS_DRA_INCONSISTENT_DIT (8443)
value ERROR_DS_DRA_INTERNAL_ERROR (8442)
value ERROR_DS_DRA_INVALID_PARAMETER (8437)
value ERROR_DS_DRA_MAIL_PROBLEM (8447)
value ERROR_DS_DRA_MISSING_KRBTGT_SECRET (8633)
value ERROR_DS_DRA_MISSING_PARENT (8460)
value ERROR_DS_DRA_NAME_COLLISION (8458)
value ERROR_DS_DRA_NOT_SUPPORTED (8454)
value ERROR_DS_DRA_NO_REPLICA (8452)
value ERROR_DS_DRA_OBJ_IS_REP_SOURCE (8450)
value ERROR_DS_DRA_OBJ_NC_MISMATCH (8545)
value ERROR_DS_DRA_OUT_OF_MEM (8446)
value ERROR_DS_DRA_OUT_SCHEDULE_WINDOW (8617)
value ERROR_DS_DRA_PREEMPTED (8461)
value ERROR_DS_DRA_RECYCLED_TARGET (8639)
value ERROR_DS_DRA_REF_ALREADY_EXISTS (8448)
value ERROR_DS_DRA_REF_NOT_FOUND (8449)
value ERROR_DS_DRA_REPL_PENDING (8477)
value ERROR_DS_DRA_RPC_CANCELLED (8455)
value ERROR_DS_DRA_SCHEMA_CONFLICT (8543)
value ERROR_DS_DRA_SCHEMA_INFO_SHIP (8542)
value ERROR_DS_DRA_SCHEMA_MISMATCH (8418)
value ERROR_DS_DRA_SECRETS_DENIED (8630)
value ERROR_DS_DRA_SHUTDOWN (8463)
value ERROR_DS_DRA_SINK_DISABLED (8457)
value ERROR_DS_DRA_SOURCE_DISABLED (8456)
value ERROR_DS_DRA_SOURCE_IS_PARTIAL_REPLICA (8465)
value ERROR_DS_DRA_SOURCE_REINSTALLED (8459)
value ERROR_DS_DRS_EXTENSIONS_CHANGED (8594)
value ERROR_DS_DSA_MUST_BE_INT_MASTER (8342)
value ERROR_DS_DST_DOMAIN_NOT_NATIVE (8496)
value ERROR_DS_DST_NC_MISMATCH (8486)
value ERROR_DS_DS_REQUIRED (8478)
value ERROR_DS_DUPLICATE_ID_FOUND (8605)
value ERROR_DS_DUP_LDAP_DISPLAY_NAME (8382)
value ERROR_DS_DUP_LINK_ID (8468)
value ERROR_DS_DUP_MAPI_ID (8380)
value ERROR_DS_DUP_MSDS_INTID (8597)
value ERROR_DS_DUP_OID (8379)
value ERROR_DS_DUP_RDN (8378)
value ERROR_DS_DUP_SCHEMA_ID_GUID (8381)
value ERROR_DS_ENCODING_ERROR (8252)
value ERROR_DS_EPOCH_MISMATCH (8483)
value ERROR_DS_EXISTING_AD_CHILD_NC (8613)
value ERROR_DS_EXISTS_IN_AUX_CLS (8393)
value ERROR_DS_EXISTS_IN_MAY_HAVE (8386)
value ERROR_DS_EXISTS_IN_MUST_HAVE (8385)
value ERROR_DS_EXISTS_IN_POSS_SUP (8395)
value ERROR_DS_EXISTS_IN_RDNATTID (8598)
value ERROR_DS_EXISTS_IN_SUB_CLS (8394)
value ERROR_DS_FILTER_UNKNOWN (8254)
value ERROR_DS_FILTER_USES_CONTRUCTED_ATTRS (8555)
value ERROR_DS_FLAT_NAME_EXISTS_IN_FOREST (8635)
value ERROR_DS_FOREST_VERSION_TOO_HIGH (8563)
value ERROR_DS_FOREST_VERSION_TOO_LOW (8565)
value ERROR_DS_GCVERIFY_ERROR (8417)
value ERROR_DS_GC_NOT_AVAILABLE (8217)
value ERROR_DS_GC_REQUIRED (8547)
value ERROR_DS_GENERIC_ERROR (8341)
value ERROR_DS_GLOBAL_CANT_HAVE_CROSSDOMAIN_MEMBER (8519)
value ERROR_DS_GLOBAL_CANT_HAVE_LOCAL_MEMBER (8516)
value ERROR_DS_GLOBAL_CANT_HAVE_UNIVERSAL_MEMBER (8517)
value ERROR_DS_GOVERNSID_MISSING (8410)
value ERROR_DS_GROUP_CONVERSION_ERROR (8607)
value ERROR_DS_HAVE_PRIMARY_MEMBERS (8521)
value ERROR_DS_HIERARCHY_TABLE_MALLOC_FAILED (8429)
value ERROR_DS_HIERARCHY_TABLE_TOO_DEEP (8628)
value ERROR_DS_HIGH_ADLDS_FFL (8641)
value ERROR_DS_HIGH_DSA_VERSION (8642)
value ERROR_DS_ILLEGAL_BASE_SCHEMA_MOD (8507)
value ERROR_DS_ILLEGAL_MOD_OPERATION (8311)
value ERROR_DS_ILLEGAL_SUPERIOR (8345)
value ERROR_DS_ILLEGAL_XDOM_MOVE_OPERATION (8492)
value ERROR_DS_INAPPROPRIATE_AUTH (8233)
value ERROR_DS_INAPPROPRIATE_MATCHING (8238)
value ERROR_DS_INCOMPATIBLE_CONTROLS_USED (8574)
value ERROR_DS_INCOMPATIBLE_VERSION (8567)
value ERROR_DS_INCORRECT_ROLE_OWNER (8210)
value ERROR_DS_INIT_FAILURE (8532)
value ERROR_DS_INIT_FAILURE_CONSOLE (8561)
value ERROR_DS_INSTALL_NO_SCH_VERSION_IN_INIFILE (8512)
value ERROR_DS_INSTALL_NO_SRC_SCH_VERSION (8511)
value ERROR_DS_INSTALL_SCHEMA_MISMATCH (8467)
value ERROR_DS_INSUFFICIENT_ATTR_TO_CREATE_OBJECT (8606)
value ERROR_DS_INSUFF_ACCESS_RIGHTS (8344)
value ERROR_DS_INTERNAL_FAILURE (8430)
value ERROR_DS_INVALID_ATTRIBUTE_SYNTAX (8203)
value ERROR_DS_INVALID_DMD (8360)
value ERROR_DS_INVALID_DN_SYNTAX (8242)
value ERROR_DS_INVALID_GROUP_TYPE (8513)
value ERROR_DS_INVALID_LDAP_DISPLAY_NAME (8479)
value ERROR_DS_INVALID_NAME_FOR_SPN (8554)
value ERROR_DS_INVALID_ROLE_OWNER (8366)
value ERROR_DS_INVALID_SCRIPT (8600)
value ERROR_DS_INVALID_SEARCH_FLAG (8500)
value ERROR_DS_INVALID_SEARCH_FLAG_SUBTREE (8626)
value ERROR_DS_INVALID_SEARCH_FLAG_TUPLE (8627)
value ERROR_DS_IS_LEAF (8243)
value ERROR_DS_KEY_NOT_UNIQUE (8527)
value ERROR_DS_LDAP_SEND_QUEUE_FULL (8616)
value ERROR_DS_LINK_ID_NOT_AVAILABLE (8577)
value ERROR_DS_LOCAL_CANT_HAVE_CROSSDOMAIN_LOCAL_MEMBER (8520)
value ERROR_DS_LOCAL_ERROR (8251)
value ERROR_DS_LOCAL_MEMBER_OF_LOCAL_ONLY (8548)
value ERROR_DS_LOOP_DETECT (8246)
value ERROR_DS_LOW_ADLDS_FFL (8643)
value ERROR_DS_LOW_DSA_VERSION (8568)
value ERROR_DS_MACHINE_ACCOUNT_QUOTA_EXCEEDED (8557)
value ERROR_DS_MAPI_ID_NOT_AVAILABLE (8632)
value ERROR_DS_MASTERDSA_REQUIRED (8314)
value ERROR_DS_MAX_OBJ_SIZE_EXCEEDED (8304)
value ERROR_DS_MEMBERSHIP_EVALUATED_LOCALLY (8201)
value ERROR_DS_MISSING_EXPECTED_ATT (8411)
value ERROR_DS_MISSING_FOREST_TRUST (8649)
value ERROR_DS_MISSING_FSMO_SETTINGS (8434)
value ERROR_DS_MISSING_INFRASTRUCTURE_CONTAINER (8497)
value ERROR_DS_MISSING_REQUIRED_ATT (8316)
value ERROR_DS_MISSING_SUPREF (8406)
value ERROR_DS_MODIFYDN_DISALLOWED_BY_FLAG (8581)
value ERROR_DS_MODIFYDN_DISALLOWED_BY_INSTANCE_TYPE (8579)
value ERROR_DS_MODIFYDN_WRONG_GRANDPARENT (8582)
value ERROR_DS_MUST_BE_RUN_ON_DST_DC (8558)
value ERROR_DS_NAME_ERROR_DOMAIN_ONLY (8473)
value ERROR_DS_NAME_ERROR_NOT_FOUND (8470)
value ERROR_DS_NAME_ERROR_NOT_UNIQUE (8471)
value ERROR_DS_NAME_ERROR_NO_MAPPING (8472)
value ERROR_DS_NAME_ERROR_NO_SYNTACTICAL_MAPPING (8474)
value ERROR_DS_NAME_ERROR_RESOLVING (8469)
value ERROR_DS_NAME_ERROR_TRUST_REFERRAL (8583)
value ERROR_DS_NAME_NOT_UNIQUE (8571)
value ERROR_DS_NAME_REFERENCE_INVALID (8373)
value ERROR_DS_NAME_TOO_LONG (8348)
value ERROR_DS_NAME_TOO_MANY_PARTS (8347)
value ERROR_DS_NAME_TYPE_UNKNOWN (8351)
value ERROR_DS_NAME_UNPARSEABLE (8350)
value ERROR_DS_NAME_VALUE_TOO_LONG (8349)
value ERROR_DS_NAMING_MASTER_GC (8523)
value ERROR_DS_NAMING_VIOLATION (8247)
value ERROR_DS_NCNAME_MISSING_CR_REF (8412)
value ERROR_DS_NCNAME_MUST_BE_NC (8357)
value ERROR_DS_NC_MUST_HAVE_NC_PARENT (8494)
value ERROR_DS_NC_STILL_HAS_DSAS (8546)
value ERROR_DS_NONEXISTENT_MAY_HAVE (8387)
value ERROR_DS_NONEXISTENT_MUST_HAVE (8388)
value ERROR_DS_NONEXISTENT_POSS_SUP (8390)
value ERROR_DS_NONSAFE_SCHEMA_CHANGE (8508)
value ERROR_DS_NON_ASQ_SEARCH (8624)
value ERROR_DS_NON_BASE_SEARCH (8480)
value ERROR_DS_NOTIFY_FILTER_TOO_COMPLEX (8377)
value ERROR_DS_NOT_AN_OBJECT (8352)
value ERROR_DS_NOT_AUTHORITIVE_FOR_DST_NC (8487)
value ERROR_DS_NOT_CLOSEST (8588)
value ERROR_DS_NOT_INSTALLED (8200)
value ERROR_DS_NOT_ON_BACKLINK (8362)
value ERROR_DS_NOT_SUPPORTED (8256)
value ERROR_DS_NOT_SUPPORTED_SORT_ORDER (8570)
value ERROR_DS_NO_ATTRIBUTE_OR_VALUE (8202)
value ERROR_DS_NO_BEHAVIOR_VERSION_IN_MIXEDDOMAIN (8569)
value ERROR_DS_NO_CHAINED_EVAL (8328)
value ERROR_DS_NO_CHAINING (8327)
value ERROR_DS_NO_CHECKPOINT_WITH_PDC (8551)
value ERROR_DS_NO_CROSSREF_FOR_NC (8363)
value ERROR_DS_NO_DELETED_NAME (8355)
value ERROR_DS_NO_FPO_IN_UNIVERSAL_GROUPS (8549)
value ERROR_DS_NO_MORE_RIDS (8209)
value ERROR_DS_NO_MSDS_INTID (8596)
value ERROR_DS_NO_NEST_GLOBALGROUP_IN_MIXEDDOMAIN (8514)
value ERROR_DS_NO_NEST_LOCALGROUP_IN_MIXEDDOMAIN (8515)
value ERROR_DS_NO_NTDSA_OBJECT (8623)
value ERROR_DS_NO_OBJECT_MOVE_IN_SCHEMA_NC (8580)
value ERROR_DS_NO_PARENT_OBJECT (8329)
value ERROR_DS_NO_PKT_PRIVACY_ON_CONNECTION (8533)
value ERROR_DS_NO_RDN_DEFINED_IN_SCHEMA (8306)
value ERROR_DS_NO_REF_DOMAIN (8575)
value ERROR_DS_NO_REQUESTED_ATTS_FOUND (8308)
value ERROR_DS_NO_RESULTS_RETURNED (8257)
value ERROR_DS_NO_RIDS_ALLOCATED (8208)
value ERROR_DS_NO_SERVER_OBJECT (8622)
value ERROR_DS_NO_SUCH_OBJECT (8240)
value ERROR_DS_NO_TREE_DELETE_ABOVE_NC (8501)
value ERROR_DS_NTDSCRIPT_PROCESS_ERROR (8592)
value ERROR_DS_NTDSCRIPT_SYNTAX_ERROR (8591)
value ERROR_DS_OBJECT_BEING_REMOVED (8339)
value ERROR_DS_OBJECT_CLASS_REQUIRED (8315)
value ERROR_DS_OBJECT_RESULTS_TOO_LARGE (8248)
value ERROR_DS_OBJ_CLASS_NOT_DEFINED (8371)
value ERROR_DS_OBJ_CLASS_NOT_SUBCLASS (8372)
value ERROR_DS_OBJ_CLASS_VIOLATION (8212)
value ERROR_DS_OBJ_GUID_EXISTS (8361)
value ERROR_DS_OBJ_NOT_FOUND (8333)
value ERROR_DS_OBJ_STRING_NAME_EXISTS (8305)
value ERROR_DS_OBJ_TOO_LARGE (8312)
value ERROR_DS_OFFSET_RANGE_ERROR (8262)
value ERROR_DS_OID_MAPPED_GROUP_CANT_HAVE_MEMBERS (8637)
value ERROR_DS_OID_NOT_FOUND (8638)
value ERROR_DS_OPERATIONS_ERROR (8224)
value ERROR_DS_OUT_OF_SCOPE (8338)
value ERROR_DS_OUT_OF_VERSION_STORE (8573)
value ERROR_DS_PARAM_ERROR (8255)
value ERROR_DS_PARENT_IS_AN_ALIAS (8330)
value ERROR_DS_PDC_OPERATION_IN_PROGRESS (8490)
value ERROR_DS_PER_ATTRIBUTE_AUTHZ_FAILED_DURING_ADD (8652)
value ERROR_DS_POLICY_NOT_KNOWN (8618)
value ERROR_DS_PROTOCOL_ERROR (8225)
value ERROR_DS_RANGE_CONSTRAINT (8322)
value ERROR_DS_RDN_DOESNT_MATCH_SCHEMA (8307)
value ERROR_DS_RECALCSCHEMA_FAILED (8396)
value ERROR_DS_REFERRAL (8235)
value ERROR_DS_REFERRAL_LIMIT_EXCEEDED (8260)
value ERROR_DS_REFUSING_FSMO_ROLES (8433)
value ERROR_DS_REMOTE_CROSSREF_OP_FAILED (8601)
value ERROR_DS_REPLICATOR_ONLY (8370)
value ERROR_DS_REPLICA_SET_CHANGE_NOT_ALLOWED_ON_DISABLED_CR (8595)
value ERROR_DS_REPL_LIFETIME_EXCEEDED (8614)
value ERROR_DS_RESERVED_LINK_ID (8576)
value ERROR_DS_RESERVED_MAPI_ID (8631)
value ERROR_DS_RIDMGR_DISABLED (8263)
value ERROR_DS_RIDMGR_INIT_ERROR (8211)
value ERROR_DS_ROLE_NOT_VERIFIED (8610)
value ERROR_DS_ROOT_CANT_BE_SUBREF (8326)
value ERROR_DS_ROOT_MUST_BE_NC (8301)
value ERROR_DS_ROOT_REQUIRES_CLASS_TOP (8432)
value ERROR_DS_SAM_INIT_FAILURE (8504)
value ERROR_DS_SAM_INIT_FAILURE_CONSOLE (8562)
value ERROR_DS_SAM_NEED_BOOTKEY_FLOPPY (8530)
value ERROR_DS_SAM_NEED_BOOTKEY_PASSWORD (8529)
value ERROR_DS_SCHEMA_ALLOC_FAILED (8415)
value ERROR_DS_SCHEMA_NOT_LOADED (8414)
value ERROR_DS_SCHEMA_UPDATE_DISALLOWED (8509)
value ERROR_DS_SECURITY_CHECKING_ERROR (8413)
value ERROR_DS_SECURITY_ILLEGAL_MODIFY (8423)
value ERROR_DS_SEC_DESC_INVALID (8354)
value ERROR_DS_SEC_DESC_TOO_SHORT (8353)
value ERROR_DS_SEMANTIC_ATT_TEST (8383)
value ERROR_DS_SENSITIVE_GROUP_VIOLATION (8505)
value ERROR_DS_SERVER_DOWN (8250)
value ERROR_DS_SHUTTING_DOWN (8364)
value ERROR_DS_SINGLE_USER_MODE_FAILED (8590)
value ERROR_DS_SINGLE_VALUE_CONSTRAINT (8321)
value ERROR_DS_SIZELIMIT_EXCEEDED (8227)
value ERROR_DS_SORT_CONTROL_MISSING (8261)
value ERROR_DS_SOURCE_AUDITING_NOT_ENABLED (8552)
value ERROR_DS_SOURCE_DOMAIN_IN_FOREST (8534)
value ERROR_DS_SPN_VALUE_NOT_UNIQUE_IN_FOREST (8647)
value ERROR_DS_SRC_AND_DST_NC_IDENTICAL (8485)
value ERROR_DS_SRC_AND_DST_OBJECT_CLASS_MISMATCH (8540)
value ERROR_DS_SRC_GUID_MISMATCH (8488)
value ERROR_DS_SRC_NAME_MISMATCH (8484)
value ERROR_DS_SRC_OBJ_NOT_GROUP_OR_USER (8538)
value ERROR_DS_SRC_SID_EXISTS_IN_FOREST (8539)
value ERROR_DS_STRING_SD_CONVERSION_FAILED (8522)
value ERROR_DS_STRONG_AUTH_REQUIRED (8232)
value ERROR_DS_SUBREF_MUST_HAVE_PARENT (8356)
value ERROR_DS_SUBTREE_NOTIFY_NOT_NC_HEAD (8376)
value ERROR_DS_SUB_CLS_TEST_FAIL (8391)
value ERROR_DS_SYNTAX_MISMATCH (8384)
value ERROR_DS_THREAD_LIMIT_EXCEEDED (8587)
value ERROR_DS_TIMELIMIT_EXCEEDED (8226)
value ERROR_DS_TREE_DELETE_NOT_FINISHED (8397)
value ERROR_DS_UNABLE_TO_SURRENDER_ROLES (8435)
value ERROR_DS_UNAVAILABLE (8207)
value ERROR_DS_UNAVAILABLE_CRIT_EXTENSION (8236)
value ERROR_DS_UNDELETE_SAM_VALIDATION_FAILED (8645)
value ERROR_DS_UNICODEPWD_NOT_IN_QUOTES (8556)
value ERROR_DS_UNIVERSAL_CANT_HAVE_LOCAL_MEMBER (8518)
value ERROR_DS_UNKNOWN_ERROR (8431)
value ERROR_DS_UNKNOWN_OPERATION (8365)
value ERROR_DS_UNWILLING_TO_PERFORM (8245)
value ERROR_DS_UPN_VALUE_NOT_UNIQUE_IN_FOREST (8648)
value ERROR_DS_USER_BUFFER_TO_SMALL (8309)
value ERROR_DS_VALUE_KEY_NOT_UNIQUE (8650)
value ERROR_DS_VERSION_CHECK_FAILURE (643)
value ERROR_DS_WKO_CONTAINER_CANNOT_BE_SPECIAL (8611)
value ERROR_DS_WRONG_LINKED_ATT_SYNTAX (8528)
value ERROR_DS_WRONG_OM_OBJ_CLASS (8476)
value ERROR_DUPLICATE_PRIVILEGES (311)
value ERROR_DUPLICATE_SERVICE_NAME (1078)
value ERROR_DUPLICATE_TAG (2014)
value ERROR_DUP_DOMAINNAME (1221)
value ERROR_DUP_NAME (52)
value ERROR_DYNAMIC_CODE_BLOCKED (1655)
value ERROR_DYNLINK_FROM_INVALID_RING (196)
value ERROR_EAS_DIDNT_FIT (275)
value ERROR_EAS_NOT_SUPPORTED (282)
value ERROR_EA_ACCESS_DENIED (994)
value ERROR_EA_FILE_CORRUPT (276)
value ERROR_EA_LIST_INCONSISTENT (255)
value ERROR_EA_TABLE_FULL (277)
value ERROR_EC_CIRCULAR_FORWARDING (15082)
value ERROR_EC_CREDSTORE_FULL (15083)
value ERROR_EC_CRED_NOT_FOUND (15084)
value ERROR_EC_LOG_DISABLED (15081)
value ERROR_EC_NO_ACTIVE_CHANNEL (15085)
value ERROR_EC_SUBSCRIPTION_CANNOT_ACTIVATE (15080)
value ERROR_EDP_DPL_POLICY_CANT_BE_SATISFIED (357)
value ERROR_EDP_POLICY_DENIES_OPERATION (356)
value ERROR_EFS_ALG_BLOB_TOO_BIG (6013)
value ERROR_EFS_DISABLED (6015)
value ERROR_EFS_NOT_ALLOWED_IN_TRANSACTION (6831)
value ERROR_EFS_SERVER_NOT_TRUSTED (6011)
value ERROR_EFS_VERSION_NOT_SUPPORT (6016)
value ERROR_ELEVATION_REQUIRED (740)
value ERROR_EMPTY (4306)
value ERROR_ENCLAVE_FAILURE (349)
value ERROR_ENCLAVE_NOT_TERMINATED (814)
value ERROR_ENCLAVE_VIOLATION (815)
value ERROR_ENCRYPTED_FILE_NOT_SUPPORTED (489)
value ERROR_ENCRYPTED_IO_NOT_POSSIBLE (808)
value ERROR_ENCRYPTING_METADATA_DISALLOWED (431)
value ERROR_ENCRYPTION_DISABLED (430)
value ERROR_ENCRYPTION_FAILED (6000)
value ERROR_ENCRYPTION_POLICY_DENIES_OPERATION (6022)
value ERROR_END_OF_MEDIA (1100)
value ERROR_ENLISTMENT_NOT_FOUND (6717)
value ERROR_ENLISTMENT_NOT_SUPERIOR (6820)
value ERROR_ENVVAR_NOT_FOUND (203)
value ERROR_EOM_OVERFLOW (1129)
value ERROR_ERRORS_ENCOUNTERED (774)
value ERROR_EVALUATION_EXPIRATION (622)
value ERROR_EVENTLOG_CANT_START (1501)
value ERROR_EVENTLOG_FILE_CHANGED (1503)
value ERROR_EVENTLOG_FILE_CORRUPT (1500)
value ERROR_EVENT_DONE (710)
value ERROR_EVENT_PENDING (711)
value ERROR_EVT_CANNOT_OPEN_CHANNEL_OF_QUERY (15036)
value ERROR_EVT_CHANNEL_CANNOT_ACTIVATE (15025)
value ERROR_EVT_CHANNEL_NOT_FOUND (15007)
value ERROR_EVT_CONFIGURATION_ERROR (15010)
value ERROR_EVT_EVENT_DEFINITION_NOT_FOUND (15032)
value ERROR_EVT_EVENT_TEMPLATE_NOT_FOUND (15003)
value ERROR_EVT_FILTER_ALREADYSCOPED (15014)
value ERROR_EVT_FILTER_INVARG (15016)
value ERROR_EVT_FILTER_INVTEST (15017)
value ERROR_EVT_FILTER_INVTYPE (15018)
value ERROR_EVT_FILTER_NOTELTSET (15015)
value ERROR_EVT_FILTER_OUT_OF_RANGE (15038)
value ERROR_EVT_FILTER_PARSEERR (15019)
value ERROR_EVT_FILTER_TOO_COMPLEX (15026)
value ERROR_EVT_FILTER_UNEXPECTEDTOKEN (15021)
value ERROR_EVT_FILTER_UNSUPPORTEDOP (15020)
value ERROR_EVT_INVALID_CHANNEL_PATH (15000)
value ERROR_EVT_INVALID_CHANNEL_PROPERTY_VALUE (15023)
value ERROR_EVT_INVALID_EVENT_DATA (15005)
value ERROR_EVT_INVALID_OPERATION_OVER_ENABLED_DIRECT_CHANNEL (15022)
value ERROR_EVT_INVALID_PUBLISHER_NAME (15004)
value ERROR_EVT_INVALID_PUBLISHER_PROPERTY_VALUE (15024)
value ERROR_EVT_INVALID_QUERY (15001)
value ERROR_EVT_MALFORMED_XML_TEXT (15008)
value ERROR_EVT_MAX_INSERTS_REACHED (15031)
value ERROR_EVT_MESSAGE_ID_NOT_FOUND (15028)
value ERROR_EVT_MESSAGE_LOCALE_NOT_FOUND (15033)
value ERROR_EVT_MESSAGE_NOT_FOUND (15027)
value ERROR_EVT_NON_VALIDATING_MSXML (15013)
value ERROR_EVT_PUBLISHER_DISABLED (15037)
value ERROR_EVT_PUBLISHER_METADATA_NOT_FOUND (15002)
value ERROR_EVT_QUERY_RESULT_INVALID_POSITION (15012)
value ERROR_EVT_QUERY_RESULT_STALE (15011)
value ERROR_EVT_SUBSCRIPTION_TO_DIRECT_CHANNEL (15009)
value ERROR_EVT_UNRESOLVED_PARAMETER_INSERT (15030)
value ERROR_EVT_UNRESOLVED_VALUE_INSERT (15029)
value ERROR_EVT_VERSION_TOO_NEW (15035)
value ERROR_EVT_VERSION_TOO_OLD (15034)
value ERROR_EXCEPTION_IN_RESOURCE_CALL (5930)
value ERROR_EXCEPTION_IN_SERVICE (1064)
value ERROR_EXCL_SEM_ALREADY_OWNED (101)
value ERROR_EXE_CANNOT_MODIFY_SIGNED_BINARY (217)
value ERROR_EXE_CANNOT_MODIFY_STRONG_SIGNED_BINARY (218)
value ERROR_EXE_MACHINE_TYPE_MISMATCH (216)
value ERROR_EXE_MARKED_INVALID (192)
value ERROR_EXPIRED_HANDLE (6854)
value ERROR_EXTENDED_ERROR (1208)
value ERROR_EXTERNAL_BACKING_PROVIDER_UNKNOWN (343)
value ERROR_EXTERNAL_SYSKEY_NOT_SUPPORTED (399)
value ERROR_EXTRANEOUS_INFORMATION (677)
value ERROR_FAILED_DRIVER_ENTRY (647)
value ERROR_FAILED_SERVICE_CONTROLLER_CONNECT (1063)
value ERROR_FAIL_FAST_EXCEPTION (1653)
value ERROR_FAIL_NOACTION_REBOOT (350)
value ERROR_FAIL_REBOOT_INITIATED (3018)
value ERROR_FAIL_REBOOT_REQUIRED (3017)
value ERROR_FAIL_RESTART (352)
value ERROR_FAIL_SHUTDOWN (351)
value ERROR_FATAL_APP_EXIT (713)
value ERROR_FILEMARK_DETECTED (1101)
value ERROR_FILENAME_EXCED_RANGE (206)
value ERROR_FILE_CHECKED_OUT (220)
value ERROR_FILE_CORRUPT (1392)
value ERROR_FILE_ENCRYPTED (6002)
value ERROR_FILE_EXISTS (80)
value ERROR_FILE_HANDLE_REVOKED (806)
value ERROR_FILE_IDENTITY_NOT_PERSISTENT (6823)
value ERROR_FILE_INVALID (1006)
value ERROR_FILE_LEVEL_TRIM_NOT_SUPPORTED (326)
value ERROR_FILE_METADATA_OPTIMIZATION_IN_PROGRESS (809)
value ERROR_FILE_NOT_ENCRYPTED (6007)
value ERROR_FILE_NOT_FOUND (2)
value ERROR_FILE_NOT_SUPPORTED (425)
value ERROR_FILE_OFFLINE (4350)
value ERROR_FILE_PROTECTED_UNDER_DPL (406)
value ERROR_FILE_READ_ONLY (6009)
value ERROR_FILE_SHARE_RESOURCE_CONFLICT (5938)
value ERROR_FILE_SNAP_INVALID_PARAMETER (440)
value ERROR_FILE_SNAP_IN_PROGRESS (435)
value ERROR_FILE_SNAP_IO_NOT_COORDINATED (438)
value ERROR_FILE_SNAP_MODIFY_NOT_SUPPORTED (437)
value ERROR_FILE_SNAP_UNEXPECTED_ERROR (439)
value ERROR_FILE_SNAP_USER_SECTION_NOT_SUPPORTED (436)
value ERROR_FILE_SYSTEM_LIMITATION (665)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_BUSY (371)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_INVALID_OPERATION (385)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_METADATA_CORRUPT (370)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_PROVIDER_UNKNOWN (372)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_UNAVAILABLE (369)
value ERROR_FILE_TOO_LARGE (223)
value ERROR_FIRMWARE_UPDATED (728)
value ERROR_FLOATED_SECTION (6846)
value ERROR_FLOAT_MULTIPLE_FAULTS (630)
value ERROR_FLOAT_MULTIPLE_TRAPS (631)
value ERROR_FLOPPY_BAD_REGISTERS (1125)
value ERROR_FLOPPY_ID_MARK_NOT_FOUND (1122)
value ERROR_FLOPPY_UNKNOWN_ERROR (1124)
value ERROR_FLOPPY_VOLUME (584)
value ERROR_FLOPPY_WRONG_CYLINDER (1123)
value ERROR_FLT_ALREADY_ENLISTED (_HRESULT_TYPEDEF_(0x801F001BL))
value ERROR_FLT_CBDQ_DISABLED (_HRESULT_TYPEDEF_(0x801F000EL))
value ERROR_FLT_CONTEXT_ALLOCATION_NOT_FOUND (_HRESULT_TYPEDEF_(0x801F0016L))
value ERROR_FLT_CONTEXT_ALREADY_DEFINED (_HRESULT_TYPEDEF_(0x801F0002L))
value ERROR_FLT_CONTEXT_ALREADY_LINKED (_HRESULT_TYPEDEF_(0x801F001CL))
value ERROR_FLT_DELETING_OBJECT (_HRESULT_TYPEDEF_(0x801F000BL))
value ERROR_FLT_DISALLOW_FAST_IO (_HRESULT_TYPEDEF_(0x801F0004L))
value ERROR_FLT_DO_NOT_ATTACH (_HRESULT_TYPEDEF_(0x801F000FL))
value ERROR_FLT_DO_NOT_DETACH (_HRESULT_TYPEDEF_(0x801F0010L))
value ERROR_FLT_DUPLICATE_ENTRY (_HRESULT_TYPEDEF_(0x801F000DL))
value ERROR_FLT_FILTER_NOT_FOUND (_HRESULT_TYPEDEF_(0x801F0013L))
value ERROR_FLT_FILTER_NOT_READY (_HRESULT_TYPEDEF_(0x801F0008L))
value ERROR_FLT_INSTANCE_ALTITUDE_COLLISION (_HRESULT_TYPEDEF_(0x801F0011L))
value ERROR_FLT_INSTANCE_NAME_COLLISION (_HRESULT_TYPEDEF_(0x801F0012L))
value ERROR_FLT_INSTANCE_NOT_FOUND (_HRESULT_TYPEDEF_(0x801F0015L))
value ERROR_FLT_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x801F000AL))
value ERROR_FLT_INVALID_ASYNCHRONOUS_REQUEST (_HRESULT_TYPEDEF_(0x801F0003L))
value ERROR_FLT_INVALID_CONTEXT_REGISTRATION (_HRESULT_TYPEDEF_(0x801F0017L))
value ERROR_FLT_INVALID_NAME_REQUEST (_HRESULT_TYPEDEF_(0x801F0005L))
value ERROR_FLT_IO_COMPLETE (_HRESULT_TYPEDEF_(0x001F0001L))
value ERROR_FLT_MUST_BE_NONPAGED_POOL (_HRESULT_TYPEDEF_(0x801F000CL))
value ERROR_FLT_NAME_CACHE_MISS (_HRESULT_TYPEDEF_(0x801F0018L))
value ERROR_FLT_NOT_INITIALIZED (_HRESULT_TYPEDEF_(0x801F0007L))
value ERROR_FLT_NOT_SAFE_TO_POST_OPERATION (_HRESULT_TYPEDEF_(0x801F0006L))
value ERROR_FLT_NO_DEVICE_OBJECT (_HRESULT_TYPEDEF_(0x801F0019L))
value ERROR_FLT_NO_HANDLER_DEFINED (_HRESULT_TYPEDEF_(0x801F0001L))
value ERROR_FLT_NO_WAITER_FOR_REPLY (_HRESULT_TYPEDEF_(0x801F0020L))
value ERROR_FLT_POST_OPERATION_CLEANUP (_HRESULT_TYPEDEF_(0x801F0009L))
value ERROR_FLT_REGISTRATION_BUSY (_HRESULT_TYPEDEF_(0x801F0023L))
value ERROR_FLT_VOLUME_ALREADY_MOUNTED (_HRESULT_TYPEDEF_(0x801F001AL))
value ERROR_FLT_VOLUME_NOT_FOUND (_HRESULT_TYPEDEF_(0x801F0014L))
value ERROR_FLT_WCOS_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x801F0024L))
value ERROR_FORMS_AUTH_REQUIRED (224)
value ERROR_FOUND_OUT_OF_SCOPE (601)
value ERROR_FSFILTER_OP_COMPLETED_SUCCESSFULLY (762)
value ERROR_FS_DRIVER_REQUIRED (588)
value ERROR_FS_METADATA_INCONSISTENT (510)
value ERROR_FT_DI_SCAN_REQUIRED (339)
value ERROR_FT_READ_FAILURE (415)
value ERROR_FT_READ_FROM_COPY_FAILURE (818)
value ERROR_FT_READ_RECOVERY_FROM_BACKUP (704)
value ERROR_FT_WRITE_FAILURE (338)
value ERROR_FT_WRITE_RECOVERY (705)
value ERROR_FULLSCREEN_MODE (1007)
value ERROR_FULL_BACKUP (4004)
value ERROR_FUNCTION_FAILED (1627)
value ERROR_FUNCTION_NOT_CALLED (1626)
value ERROR_GDI_HANDLE_LEAK (373)
value ERROR_GENERIC_COMMAND_FAILED (14109)
value ERROR_GENERIC_NOT_MAPPED (1360)
value ERROR_GEN_FAILURE (31)
value ERROR_GLOBAL_ONLY_HOOK (1429)
value ERROR_GPIO_CLIENT_INFORMATION_INVALID (15322)
value ERROR_GPIO_INCOMPATIBLE_CONNECT_MODE (15326)
value ERROR_GPIO_INTERRUPT_ALREADY_UNMASKED (15327)
value ERROR_GPIO_INVALID_REGISTRATION_PACKET (15324)
value ERROR_GPIO_OPERATION_DENIED (15325)
value ERROR_GPIO_VERSION_NOT_SUPPORTED (15323)
value ERROR_GRACEFUL_DISCONNECT (1226)
value ERROR_GRAPHICS_ADAPTER_ACCESS_NOT_EXCLUDED (_HRESULT_TYPEDEF_(0xC026243BL))
value ERROR_GRAPHICS_ADAPTER_CHAIN_NOT_READY (_HRESULT_TYPEDEF_(0xC0262433L))
value ERROR_GRAPHICS_ADAPTER_MUST_HAVE_AT_LEAST_ONE_SOURCE (_HRESULT_TYPEDEF_(0xC0262328L))
value ERROR_GRAPHICS_ADAPTER_MUST_HAVE_AT_LEAST_ONE_TARGET (_HRESULT_TYPEDEF_(0xC0262329L))
value ERROR_GRAPHICS_ADAPTER_WAS_RESET (_HRESULT_TYPEDEF_(0xC0262003L))
value ERROR_GRAPHICS_ALLOCATION_BUSY (_HRESULT_TYPEDEF_(0xC0262102L))
value ERROR_GRAPHICS_ALLOCATION_CLOSED (_HRESULT_TYPEDEF_(0xC0262112L))
value ERROR_GRAPHICS_ALLOCATION_CONTENT_LOST (_HRESULT_TYPEDEF_(0xC0262116L))
value ERROR_GRAPHICS_ALLOCATION_INVALID (_HRESULT_TYPEDEF_(0xC0262106L))
value ERROR_GRAPHICS_CANCEL_VIDPN_TOPOLOGY_AUGMENTATION (_HRESULT_TYPEDEF_(0xC026235AL))
value ERROR_GRAPHICS_CANNOTCOLORCONVERT (_HRESULT_TYPEDEF_(0xC0262008L))
value ERROR_GRAPHICS_CANT_ACCESS_ACTIVE_VIDPN (_HRESULT_TYPEDEF_(0xC0262343L))
value ERROR_GRAPHICS_CANT_EVICT_PINNED_ALLOCATION (_HRESULT_TYPEDEF_(0xC0262109L))
value ERROR_GRAPHICS_CANT_LOCK_MEMORY (_HRESULT_TYPEDEF_(0xC0262101L))
value ERROR_GRAPHICS_CANT_RENDER_LOCKED_ALLOCATION (_HRESULT_TYPEDEF_(0xC0262111L))
value ERROR_GRAPHICS_CHAINLINKS_NOT_ENUMERATED (_HRESULT_TYPEDEF_(0xC0262432L))
value ERROR_GRAPHICS_CHAINLINKS_NOT_POWERED_ON (_HRESULT_TYPEDEF_(0xC0262435L))
value ERROR_GRAPHICS_CHAINLINKS_NOT_STARTED (_HRESULT_TYPEDEF_(0xC0262434L))
value ERROR_GRAPHICS_CHILD_DESCRIPTOR_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262401L))
value ERROR_GRAPHICS_CLIENTVIDPN_NOT_SET (_HRESULT_TYPEDEF_(0xC026235CL))
value ERROR_GRAPHICS_COPP_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262501L))
value ERROR_GRAPHICS_DATASET_IS_EMPTY (_HRESULT_TYPEDEF_(0x0026234BL))
value ERROR_GRAPHICS_DDCCI_CURRENT_CURRENT_VALUE_GREATER_THAN_MAXIMUM_VALUE (_HRESULT_TYPEDEF_(0xC02625D8L))
value ERROR_GRAPHICS_DDCCI_INVALID_DATA (_HRESULT_TYPEDEF_(0xC0262585L))
value ERROR_GRAPHICS_DDCCI_INVALID_MESSAGE_CHECKSUM (_HRESULT_TYPEDEF_(0xC026258BL))
value ERROR_GRAPHICS_DDCCI_INVALID_MESSAGE_COMMAND (_HRESULT_TYPEDEF_(0xC0262589L))
value ERROR_GRAPHICS_DDCCI_INVALID_MESSAGE_LENGTH (_HRESULT_TYPEDEF_(0xC026258AL))
value ERROR_GRAPHICS_DDCCI_MONITOR_RETURNED_INVALID_TIMING_STATUS_BYTE (_HRESULT_TYPEDEF_(0xC0262586L))
value ERROR_GRAPHICS_DDCCI_VCP_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262584L))
value ERROR_GRAPHICS_DEPENDABLE_CHILD_STATUS (_HRESULT_TYPEDEF_(0x4026243CL))
value ERROR_GRAPHICS_DISPLAY_DEVICE_NOT_ATTACHED_TO_DESKTOP (_HRESULT_TYPEDEF_(0xC02625E2L))
value ERROR_GRAPHICS_DRIVER_MISMATCH (_HRESULT_TYPEDEF_(0xC0262009L))
value ERROR_GRAPHICS_EMPTY_ADAPTER_MONITOR_MODE_SUPPORT_INTERSECTION (_HRESULT_TYPEDEF_(0xC0262325L))
value ERROR_GRAPHICS_FREQUENCYRANGE_ALREADY_IN_SET (_HRESULT_TYPEDEF_(0xC026231FL))
value ERROR_GRAPHICS_FREQUENCYRANGE_NOT_IN_SET (_HRESULT_TYPEDEF_(0xC026231DL))
value ERROR_GRAPHICS_GAMMA_RAMP_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262348L))
value ERROR_GRAPHICS_GPU_EXCEPTION_ON_DEVICE (_HRESULT_TYPEDEF_(0xC0262200L))
value ERROR_GRAPHICS_INCOMPATIBLE_PRIVATE_FORMAT (_HRESULT_TYPEDEF_(0xC0262355L))
value ERROR_GRAPHICS_INCONSISTENT_DEVICE_LINK_STATE (_HRESULT_TYPEDEF_(0xC0262436L))
value ERROR_GRAPHICS_INDIRECT_DISPLAY_ABANDON_SWAPCHAIN (_HRESULT_TYPEDEF_(0xC0262012L))
value ERROR_GRAPHICS_INDIRECT_DISPLAY_DEVICE_STOPPED (_HRESULT_TYPEDEF_(0xC0262013L))
value ERROR_GRAPHICS_INSUFFICIENT_DMA_BUFFER (_HRESULT_TYPEDEF_(0xC0262001L))
value ERROR_GRAPHICS_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0xC02625E7L))
value ERROR_GRAPHICS_INVALID_ACTIVE_REGION (_HRESULT_TYPEDEF_(0xC026230BL))
value ERROR_GRAPHICS_INVALID_ALLOCATION_HANDLE (_HRESULT_TYPEDEF_(0xC0262114L))
value ERROR_GRAPHICS_INVALID_ALLOCATION_INSTANCE (_HRESULT_TYPEDEF_(0xC0262113L))
value ERROR_GRAPHICS_INVALID_ALLOCATION_USAGE (_HRESULT_TYPEDEF_(0xC0262110L))
value ERROR_GRAPHICS_INVALID_CLIENT_TYPE (_HRESULT_TYPEDEF_(0xC026235BL))
value ERROR_GRAPHICS_INVALID_COLORBASIS (_HRESULT_TYPEDEF_(0xC026233EL))
value ERROR_GRAPHICS_INVALID_COPYPROTECTION_TYPE (_HRESULT_TYPEDEF_(0xC026234FL))
value ERROR_GRAPHICS_INVALID_DISPLAY_ADAPTER (_HRESULT_TYPEDEF_(0xC0262002L))
value ERROR_GRAPHICS_INVALID_DRIVER_MODEL (_HRESULT_TYPEDEF_(0xC0262004L))
value ERROR_GRAPHICS_INVALID_FREQUENCY (_HRESULT_TYPEDEF_(0xC026230AL))
value ERROR_GRAPHICS_INVALID_GAMMA_RAMP (_HRESULT_TYPEDEF_(0xC0262347L))
value ERROR_GRAPHICS_INVALID_MODE_PRUNING_ALGORITHM (_HRESULT_TYPEDEF_(0xC0262356L))
value ERROR_GRAPHICS_INVALID_MONITORDESCRIPTOR (_HRESULT_TYPEDEF_(0xC026232BL))
value ERROR_GRAPHICS_INVALID_MONITORDESCRIPTORSET (_HRESULT_TYPEDEF_(0xC026232AL))
value ERROR_GRAPHICS_INVALID_MONITOR_CAPABILITY_ORIGIN (_HRESULT_TYPEDEF_(0xC0262357L))
value ERROR_GRAPHICS_INVALID_MONITOR_FREQUENCYRANGE (_HRESULT_TYPEDEF_(0xC026231CL))
value ERROR_GRAPHICS_INVALID_MONITOR_FREQUENCYRANGESET (_HRESULT_TYPEDEF_(0xC026231BL))
value ERROR_GRAPHICS_INVALID_MONITOR_FREQUENCYRANGE_CONSTRAINT (_HRESULT_TYPEDEF_(0xC0262358L))
value ERROR_GRAPHICS_INVALID_MONITOR_SOURCEMODESET (_HRESULT_TYPEDEF_(0xC0262321L))
value ERROR_GRAPHICS_INVALID_MONITOR_SOURCE_MODE (_HRESULT_TYPEDEF_(0xC0262322L))
value ERROR_GRAPHICS_INVALID_PATH_CONTENT_GEOMETRY_TRANSFORMATION (_HRESULT_TYPEDEF_(0xC0262345L))
value ERROR_GRAPHICS_INVALID_PATH_CONTENT_TYPE (_HRESULT_TYPEDEF_(0xC026234EL))
value ERROR_GRAPHICS_INVALID_PATH_IMPORTANCE_ORDINAL (_HRESULT_TYPEDEF_(0xC0262344L))
value ERROR_GRAPHICS_INVALID_PHYSICAL_MONITOR_HANDLE (_HRESULT_TYPEDEF_(0xC026258CL))
value ERROR_GRAPHICS_INVALID_PIXELFORMAT (_HRESULT_TYPEDEF_(0xC026233DL))
value ERROR_GRAPHICS_INVALID_PIXELVALUEACCESSMODE (_HRESULT_TYPEDEF_(0xC026233FL))
value ERROR_GRAPHICS_INVALID_POINTER (_HRESULT_TYPEDEF_(0xC02625E4L))
value ERROR_GRAPHICS_INVALID_PRIMARYSURFACE_SIZE (_HRESULT_TYPEDEF_(0xC026233AL))
value ERROR_GRAPHICS_INVALID_SCANLINE_ORDERING (_HRESULT_TYPEDEF_(0xC0262352L))
value ERROR_GRAPHICS_INVALID_STRIDE (_HRESULT_TYPEDEF_(0xC026233CL))
value ERROR_GRAPHICS_INVALID_TOTAL_REGION (_HRESULT_TYPEDEF_(0xC026230CL))
value ERROR_GRAPHICS_INVALID_VIDEOPRESENTSOURCESET (_HRESULT_TYPEDEF_(0xC0262315L))
value ERROR_GRAPHICS_INVALID_VIDEOPRESENTTARGETSET (_HRESULT_TYPEDEF_(0xC0262316L))
value ERROR_GRAPHICS_INVALID_VIDEO_PRESENT_SOURCE (_HRESULT_TYPEDEF_(0xC0262304L))
value ERROR_GRAPHICS_INVALID_VIDEO_PRESENT_SOURCE_MODE (_HRESULT_TYPEDEF_(0xC0262310L))
value ERROR_GRAPHICS_INVALID_VIDEO_PRESENT_TARGET (_HRESULT_TYPEDEF_(0xC0262305L))
value ERROR_GRAPHICS_INVALID_VIDEO_PRESENT_TARGET_MODE (_HRESULT_TYPEDEF_(0xC0262311L))
value ERROR_GRAPHICS_INVALID_VIDPN (_HRESULT_TYPEDEF_(0xC0262303L))
value ERROR_GRAPHICS_INVALID_VIDPN_PRESENT_PATH (_HRESULT_TYPEDEF_(0xC0262319L))
value ERROR_GRAPHICS_INVALID_VIDPN_SOURCEMODESET (_HRESULT_TYPEDEF_(0xC0262308L))
value ERROR_GRAPHICS_INVALID_VIDPN_TARGETMODESET (_HRESULT_TYPEDEF_(0xC0262309L))
value ERROR_GRAPHICS_INVALID_VIDPN_TARGET_SUBSET_TYPE (_HRESULT_TYPEDEF_(0xC026232FL))
value ERROR_GRAPHICS_INVALID_VIDPN_TOPOLOGY (_HRESULT_TYPEDEF_(0xC0262300L))
value ERROR_GRAPHICS_INVALID_VIDPN_TOPOLOGY_RECOMMENDATION_REASON (_HRESULT_TYPEDEF_(0xC026234DL))
value ERROR_GRAPHICS_INVALID_VISIBLEREGION_SIZE (_HRESULT_TYPEDEF_(0xC026233BL))
value ERROR_GRAPHICS_LEADLINK_NOT_ENUMERATED (_HRESULT_TYPEDEF_(0xC0262431L))
value ERROR_GRAPHICS_LEADLINK_START_DEFERRED (_HRESULT_TYPEDEF_(0x40262437L))
value ERROR_GRAPHICS_LINK_CONFIGURATION_IN_PROGRESS (_HRESULT_TYPEDEF_(0xC0262017L))
value ERROR_GRAPHICS_MAX_NUM_PATHS_REACHED (_HRESULT_TYPEDEF_(0xC0262359L))
value ERROR_GRAPHICS_MCA_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0xC0262588L))
value ERROR_GRAPHICS_MCA_INVALID_CAPABILITIES_STRING (_HRESULT_TYPEDEF_(0xC0262587L))
value ERROR_GRAPHICS_MCA_INVALID_TECHNOLOGY_TYPE_RETURNED (_HRESULT_TYPEDEF_(0xC02625DEL))
value ERROR_GRAPHICS_MCA_INVALID_VCP_VERSION (_HRESULT_TYPEDEF_(0xC02625D9L))
value ERROR_GRAPHICS_MCA_MCCS_VERSION_MISMATCH (_HRESULT_TYPEDEF_(0xC02625DBL))
value ERROR_GRAPHICS_MCA_MONITOR_VIOLATES_MCCS_SPECIFICATION (_HRESULT_TYPEDEF_(0xC02625DAL))
value ERROR_GRAPHICS_MCA_UNSUPPORTED_COLOR_TEMPERATURE (_HRESULT_TYPEDEF_(0xC02625DFL))
value ERROR_GRAPHICS_MCA_UNSUPPORTED_MCCS_VERSION (_HRESULT_TYPEDEF_(0xC02625DCL))
value ERROR_GRAPHICS_MIRRORING_DEVICES_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC02625E3L))
value ERROR_GRAPHICS_MODE_ALREADY_IN_MODESET (_HRESULT_TYPEDEF_(0xC0262314L))
value ERROR_GRAPHICS_MODE_ID_MUST_BE_UNIQUE (_HRESULT_TYPEDEF_(0xC0262324L))
value ERROR_GRAPHICS_MODE_NOT_IN_MODESET (_HRESULT_TYPEDEF_(0xC026234AL))
value ERROR_GRAPHICS_MODE_NOT_PINNED (_HRESULT_TYPEDEF_(0x00262307L))
value ERROR_GRAPHICS_MONITORDESCRIPTOR_ALREADY_IN_SET (_HRESULT_TYPEDEF_(0xC026232DL))
value ERROR_GRAPHICS_MONITORDESCRIPTOR_ID_MUST_BE_UNIQUE (_HRESULT_TYPEDEF_(0xC026232EL))
value ERROR_GRAPHICS_MONITORDESCRIPTOR_NOT_IN_SET (_HRESULT_TYPEDEF_(0xC026232CL))
value ERROR_GRAPHICS_MONITOR_COULD_NOT_BE_ASSOCIATED_WITH_ADAPTER (_HRESULT_TYPEDEF_(0xC0262334L))
value ERROR_GRAPHICS_MONITOR_NOT_CONNECTED (_HRESULT_TYPEDEF_(0xC0262338L))
value ERROR_GRAPHICS_MONITOR_NO_LONGER_EXISTS (_HRESULT_TYPEDEF_(0xC026258DL))
value ERROR_GRAPHICS_MPO_ALLOCATION_UNPINNED (_HRESULT_TYPEDEF_(0xC0262018L))
value ERROR_GRAPHICS_MULTISAMPLING_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262349L))
value ERROR_GRAPHICS_NOT_A_LINKED_ADAPTER (_HRESULT_TYPEDEF_(0xC0262430L))
value ERROR_GRAPHICS_NOT_EXCLUSIVE_MODE_OWNER (_HRESULT_TYPEDEF_(0xC0262000L))
value ERROR_GRAPHICS_NOT_POST_DEVICE_DRIVER (_HRESULT_TYPEDEF_(0xC0262438L))
value ERROR_GRAPHICS_NO_ACTIVE_VIDPN (_HRESULT_TYPEDEF_(0xC0262336L))
value ERROR_GRAPHICS_NO_AVAILABLE_IMPORTANCE_ORDINALS (_HRESULT_TYPEDEF_(0xC0262354L))
value ERROR_GRAPHICS_NO_AVAILABLE_VIDPN_TARGET (_HRESULT_TYPEDEF_(0xC0262333L))
value ERROR_GRAPHICS_NO_DISPLAY_DEVICE_CORRESPONDS_TO_NAME (_HRESULT_TYPEDEF_(0xC02625E1L))
value ERROR_GRAPHICS_NO_DISPLAY_MODE_MANAGEMENT_SUPPORT (_HRESULT_TYPEDEF_(0xC0262341L))
value ERROR_GRAPHICS_NO_MONITORS_CORRESPOND_TO_DISPLAY_DEVICE (_HRESULT_TYPEDEF_(0xC02625E5L))
value ERROR_GRAPHICS_NO_MORE_ELEMENTS_IN_DATASET (_HRESULT_TYPEDEF_(0x0026234CL))
value ERROR_GRAPHICS_NO_PREFERRED_MODE (_HRESULT_TYPEDEF_(0x0026231EL))
value ERROR_GRAPHICS_NO_RECOMMENDED_FUNCTIONAL_VIDPN (_HRESULT_TYPEDEF_(0xC0262323L))
value ERROR_GRAPHICS_NO_RECOMMENDED_VIDPN_TOPOLOGY (_HRESULT_TYPEDEF_(0xC026231AL))
value ERROR_GRAPHICS_NO_VIDEO_MEMORY (_HRESULT_TYPEDEF_(0xC0262100L))
value ERROR_GRAPHICS_NO_VIDPNMGR (_HRESULT_TYPEDEF_(0xC0262335L))
value ERROR_GRAPHICS_ONLY_CONSOLE_SESSION_SUPPORTED (_HRESULT_TYPEDEF_(0xC02625E0L))
value ERROR_GRAPHICS_OPM_ALL_HDCP_HARDWARE_ALREADY_IN_USE (_HRESULT_TYPEDEF_(0xC0262518L))
value ERROR_GRAPHICS_OPM_DRIVER_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0xC026251EL))
value ERROR_GRAPHICS_OPM_HDCP_SRM_NEVER_SET (_HRESULT_TYPEDEF_(0xC0262516L))
value ERROR_GRAPHICS_OPM_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0xC026250BL))
value ERROR_GRAPHICS_OPM_INVALID_CONFIGURATION_REQUEST (_HRESULT_TYPEDEF_(0xC0262521L))
value ERROR_GRAPHICS_OPM_INVALID_ENCRYPTED_PARAMETERS (_HRESULT_TYPEDEF_(0xC0262503L))
value ERROR_GRAPHICS_OPM_INVALID_HANDLE (_HRESULT_TYPEDEF_(0xC026250CL))
value ERROR_GRAPHICS_OPM_INVALID_INFORMATION_REQUEST (_HRESULT_TYPEDEF_(0xC026251DL))
value ERROR_GRAPHICS_OPM_INVALID_SRM (_HRESULT_TYPEDEF_(0xC0262512L))
value ERROR_GRAPHICS_OPM_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262500L))
value ERROR_GRAPHICS_OPM_NO_VIDEO_OUTPUTS_EXIST (_HRESULT_TYPEDEF_(0xC0262505L))
value ERROR_GRAPHICS_OPM_OUTPUT_DOES_NOT_SUPPORT_ACP (_HRESULT_TYPEDEF_(0xC0262514L))
value ERROR_GRAPHICS_OPM_OUTPUT_DOES_NOT_SUPPORT_CGMSA (_HRESULT_TYPEDEF_(0xC0262515L))
value ERROR_GRAPHICS_OPM_OUTPUT_DOES_NOT_SUPPORT_HDCP (_HRESULT_TYPEDEF_(0xC0262513L))
value ERROR_GRAPHICS_OPM_RESOLUTION_TOO_HIGH (_HRESULT_TYPEDEF_(0xC0262517L))
value ERROR_GRAPHICS_OPM_SESSION_TYPE_CHANGE_IN_PROGRESS (_HRESULT_TYPEDEF_(0xC026251BL))
value ERROR_GRAPHICS_OPM_SIGNALING_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262520L))
value ERROR_GRAPHICS_OPM_SPANNING_MODE_ENABLED (_HRESULT_TYPEDEF_(0xC026250FL))
value ERROR_GRAPHICS_OPM_THEATER_MODE_ENABLED (_HRESULT_TYPEDEF_(0xC0262510L))
value ERROR_GRAPHICS_OPM_VIDEO_OUTPUT_DOES_NOT_HAVE_COPP_SEMANTICS (_HRESULT_TYPEDEF_(0xC026251CL))
value ERROR_GRAPHICS_OPM_VIDEO_OUTPUT_DOES_NOT_HAVE_OPM_SEMANTICS (_HRESULT_TYPEDEF_(0xC026251FL))
value ERROR_GRAPHICS_OPM_VIDEO_OUTPUT_NO_LONGER_EXISTS (_HRESULT_TYPEDEF_(0xC026251AL))
value ERROR_GRAPHICS_PARAMETER_ARRAY_TOO_SMALL (_HRESULT_TYPEDEF_(0xC02625E6L))
value ERROR_GRAPHICS_PARTIAL_DATA_POPULATED (_HRESULT_TYPEDEF_(0x4026200AL))
value ERROR_GRAPHICS_PATH_ALREADY_IN_TOPOLOGY (_HRESULT_TYPEDEF_(0xC0262313L))
value ERROR_GRAPHICS_PATH_CONTENT_GEOMETRY_TRANSFORMATION_NOT_PINNED (_HRESULT_TYPEDEF_(0x00262351L))
value ERROR_GRAPHICS_PATH_CONTENT_GEOMETRY_TRANSFORMATION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262346L))
value ERROR_GRAPHICS_PATH_NOT_IN_TOPOLOGY (_HRESULT_TYPEDEF_(0xC0262327L))
value ERROR_GRAPHICS_PINNED_MODE_MUST_REMAIN_IN_SET (_HRESULT_TYPEDEF_(0xC0262312L))
value ERROR_GRAPHICS_POLLING_TOO_FREQUENTLY (_HRESULT_TYPEDEF_(0x40262439L))
value ERROR_GRAPHICS_PRESENT_BUFFER_NOT_BOUND (_HRESULT_TYPEDEF_(0xC0262010L))
value ERROR_GRAPHICS_PRESENT_DENIED (_HRESULT_TYPEDEF_(0xC0262007L))
value ERROR_GRAPHICS_PRESENT_INVALID_WINDOW (_HRESULT_TYPEDEF_(0xC026200FL))
value ERROR_GRAPHICS_PRESENT_MODE_CHANGED (_HRESULT_TYPEDEF_(0xC0262005L))
value ERROR_GRAPHICS_PRESENT_OCCLUDED (_HRESULT_TYPEDEF_(0xC0262006L))
value ERROR_GRAPHICS_PRESENT_REDIRECTION_DISABLED (_HRESULT_TYPEDEF_(0xC026200BL))
value ERROR_GRAPHICS_PRESENT_UNOCCLUDED (_HRESULT_TYPEDEF_(0xC026200CL))
value ERROR_GRAPHICS_PVP_HFS_FAILED (_HRESULT_TYPEDEF_(0xC0262511L))
value ERROR_GRAPHICS_PVP_INVALID_CERTIFICATE_LENGTH (_HRESULT_TYPEDEF_(0xC026250EL))
value ERROR_GRAPHICS_RESOURCES_NOT_RELATED (_HRESULT_TYPEDEF_(0xC0262330L))
value ERROR_GRAPHICS_SESSION_TYPE_CHANGE_IN_PROGRESS (_HRESULT_TYPEDEF_(0xC02605E8L))
value ERROR_GRAPHICS_SKIP_ALLOCATION_PREPARATION (_HRESULT_TYPEDEF_(0x40262201L))
value ERROR_GRAPHICS_SOURCE_ALREADY_IN_SET (_HRESULT_TYPEDEF_(0xC0262317L))
value ERROR_GRAPHICS_SOURCE_ID_MUST_BE_UNIQUE (_HRESULT_TYPEDEF_(0xC0262331L))
value ERROR_GRAPHICS_SOURCE_NOT_IN_TOPOLOGY (_HRESULT_TYPEDEF_(0xC0262339L))
value ERROR_GRAPHICS_SPECIFIED_CHILD_ALREADY_CONNECTED (_HRESULT_TYPEDEF_(0xC0262400L))
value ERROR_GRAPHICS_STALE_MODESET (_HRESULT_TYPEDEF_(0xC0262320L))
value ERROR_GRAPHICS_STALE_VIDPN_TOPOLOGY (_HRESULT_TYPEDEF_(0xC0262337L))
value ERROR_GRAPHICS_START_DEFERRED (_HRESULT_TYPEDEF_(0x4026243AL))
value ERROR_GRAPHICS_TARGET_ALREADY_IN_SET (_HRESULT_TYPEDEF_(0xC0262318L))
value ERROR_GRAPHICS_TARGET_ID_MUST_BE_UNIQUE (_HRESULT_TYPEDEF_(0xC0262332L))
value ERROR_GRAPHICS_TARGET_NOT_IN_TOPOLOGY (_HRESULT_TYPEDEF_(0xC0262340L))
value ERROR_GRAPHICS_TOO_MANY_REFERENCES (_HRESULT_TYPEDEF_(0xC0262103L))
value ERROR_GRAPHICS_TOPOLOGY_CHANGES_NOT_ALLOWED (_HRESULT_TYPEDEF_(0xC0262353L))
value ERROR_GRAPHICS_TRY_AGAIN_LATER (_HRESULT_TYPEDEF_(0xC0262104L))
value ERROR_GRAPHICS_TRY_AGAIN_NOW (_HRESULT_TYPEDEF_(0xC0262105L))
value ERROR_GRAPHICS_UAB_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262502L))
value ERROR_GRAPHICS_UNASSIGNED_MODESET_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0xC0262350L))
value ERROR_GRAPHICS_UNKNOWN_CHILD_STATUS (_HRESULT_TYPEDEF_(0x4026242FL))
value ERROR_GRAPHICS_UNSWIZZLING_APERTURE_UNAVAILABLE (_HRESULT_TYPEDEF_(0xC0262107L))
value ERROR_GRAPHICS_UNSWIZZLING_APERTURE_UNSUPPORTED (_HRESULT_TYPEDEF_(0xC0262108L))
value ERROR_GRAPHICS_VAIL_FAILED_TO_SEND_COMPOSITION_WINDOW_DPI_MESSAGE (_HRESULT_TYPEDEF_(0xC0262016L))
value ERROR_GRAPHICS_VAIL_FAILED_TO_SEND_CREATE_SUPERWETINK_MESSAGE (_HRESULT_TYPEDEF_(0xC0262014L))
value ERROR_GRAPHICS_VAIL_FAILED_TO_SEND_DESTROY_SUPERWETINK_MESSAGE (_HRESULT_TYPEDEF_(0xC0262015L))
value ERROR_GRAPHICS_VAIL_STATE_CHANGED (_HRESULT_TYPEDEF_(0xC0262011L))
value ERROR_GRAPHICS_VIDEO_PRESENT_TARGETS_LESS_THAN_SOURCES (_HRESULT_TYPEDEF_(0xC0262326L))
value ERROR_GRAPHICS_VIDPN_MODALITY_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262306L))
value ERROR_GRAPHICS_VIDPN_SOURCE_IN_USE (_HRESULT_TYPEDEF_(0xC0262342L))
value ERROR_GRAPHICS_VIDPN_TOPOLOGY_CURRENTLY_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262302L))
value ERROR_GRAPHICS_VIDPN_TOPOLOGY_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0262301L))
value ERROR_GRAPHICS_WINDOWDC_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0xC026200DL))
value ERROR_GRAPHICS_WINDOWLESS_PRESENT_DISABLED (_HRESULT_TYPEDEF_(0xC026200EL))
value ERROR_GRAPHICS_WRONG_ALLOCATION_DEVICE (_HRESULT_TYPEDEF_(0xC0262115L))
value ERROR_GROUPSET_CANT_PROVIDE (5993)
value ERROR_GROUPSET_NOT_AVAILABLE (5991)
value ERROR_GROUPSET_NOT_FOUND (5992)
value ERROR_GROUP_EXISTS (1318)
value ERROR_GROUP_NOT_AVAILABLE (5012)
value ERROR_GROUP_NOT_FOUND (5013)
value ERROR_GROUP_NOT_ONLINE (5014)
value ERROR_GUID_SUBSTITUTION_MADE (680)
value ERROR_HANDLES_CLOSED (676)
value ERROR_HANDLE_DISK_FULL (39)
value ERROR_HANDLE_EOF (38)
value ERROR_HANDLE_NO_LONGER_VALID (6815)
value ERROR_HANDLE_REVOKED (811)
value ERROR_HASH_NOT_PRESENT (15301)
value ERROR_HASH_NOT_SUPPORTED (15300)
value ERROR_HAS_SYSTEM_CRITICAL_FILES (488)
value ERROR_HEURISTIC_DAMAGE_POSSIBLE (6731)
value ERROR_HIBERNATED (726)
value ERROR_HIBERNATION_FAILURE (656)
value ERROR_HISTORY_DIRECTORY_ENTRY_DEFAULT_COUNT (8)
value ERROR_HOOK_NEEDS_HMOD (1428)
value ERROR_HOOK_NOT_INSTALLED (1431)
value ERROR_HOOK_TYPE_NOT_ALLOWED (1458)
value ERROR_HOST_DOWN (1256)
value ERROR_HOST_NODE_NOT_AVAILABLE (5005)
value ERROR_HOST_NODE_NOT_GROUP_OWNER (5016)
value ERROR_HOST_NODE_NOT_RESOURCE_OWNER (5015)
value ERROR_HOST_UNREACHABLE (1232)
value ERROR_HOTKEY_ALREADY_REGISTERED (1409)
value ERROR_HOTKEY_NOT_REGISTERED (1419)
value ERROR_HUNG_DISPLAY_DRIVER_THREAD (_HRESULT_TYPEDEF_(0x80260001L))
value ERROR_HV_ACCESS_DENIED (_NDIS_ERROR_TYPEDEF_(0xC0350006L))
value ERROR_HV_ACKNOWLEDGED (_NDIS_ERROR_TYPEDEF_(0xC0350016L))
value ERROR_HV_CPUID_FEATURE_VALIDATION (_NDIS_ERROR_TYPEDEF_(0xC035003CL))
value ERROR_HV_CPUID_XSAVE_FEATURE_VALIDATION (_NDIS_ERROR_TYPEDEF_(0xC035003DL))
value ERROR_HV_DEVICE_NOT_IN_DOMAIN (_NDIS_ERROR_TYPEDEF_(0xC0350076L))
value ERROR_HV_EVENT_BUFFER_ALREADY_FREED (_NDIS_ERROR_TYPEDEF_(0xC0350074L))
value ERROR_HV_FEATURE_UNAVAILABLE (_NDIS_ERROR_TYPEDEF_(0xC035001EL))
value ERROR_HV_INACTIVE (_NDIS_ERROR_TYPEDEF_(0xC035001CL))
value ERROR_HV_INSUFFICIENT_BUFFER (_NDIS_ERROR_TYPEDEF_(0xC0350033L))
value ERROR_HV_INSUFFICIENT_BUFFERS (_NDIS_ERROR_TYPEDEF_(0xC0350013L))
value ERROR_HV_INSUFFICIENT_CONTIGUOUS_MEMORY (_NDIS_ERROR_TYPEDEF_(0xC0350075L))
value ERROR_HV_INSUFFICIENT_CONTIGUOUS_MEMORY_MIRRORING (_NDIS_ERROR_TYPEDEF_(0xC0350082L))
value ERROR_HV_INSUFFICIENT_CONTIGUOUS_ROOT_MEMORY (_NDIS_ERROR_TYPEDEF_(0xC0350083L))
value ERROR_HV_INSUFFICIENT_CONTIGUOUS_ROOT_MEMORY_MIRRORING (_NDIS_ERROR_TYPEDEF_(0xC0350085L))
value ERROR_HV_INSUFFICIENT_DEVICE_DOMAINS (_NDIS_ERROR_TYPEDEF_(0xC0350038L))
value ERROR_HV_INSUFFICIENT_MEMORY (_NDIS_ERROR_TYPEDEF_(0xC035000BL))
value ERROR_HV_INSUFFICIENT_MEMORY_MIRRORING (_NDIS_ERROR_TYPEDEF_(0xC0350081L))
value ERROR_HV_INSUFFICIENT_ROOT_MEMORY (_NDIS_ERROR_TYPEDEF_(0xC0350073L))
value ERROR_HV_INSUFFICIENT_ROOT_MEMORY_MIRRORING (_NDIS_ERROR_TYPEDEF_(0xC0350084L))
value ERROR_HV_INVALID_ALIGNMENT (_NDIS_ERROR_TYPEDEF_(0xC0350004L))
value ERROR_HV_INVALID_CONNECTION_ID (_NDIS_ERROR_TYPEDEF_(0xC0350012L))
value ERROR_HV_INVALID_CPU_GROUP_ID (_NDIS_ERROR_TYPEDEF_(0xC035006FL))
value ERROR_HV_INVALID_CPU_GROUP_STATE (_NDIS_ERROR_TYPEDEF_(0xC0350070L))
value ERROR_HV_INVALID_DEVICE_ID (_NDIS_ERROR_TYPEDEF_(0xC0350057L))
value ERROR_HV_INVALID_DEVICE_STATE (_NDIS_ERROR_TYPEDEF_(0xC0350058L))
value ERROR_HV_INVALID_HYPERCALL_CODE (_NDIS_ERROR_TYPEDEF_(0xC0350002L))
value ERROR_HV_INVALID_HYPERCALL_INPUT (_NDIS_ERROR_TYPEDEF_(0xC0350003L))
value ERROR_HV_INVALID_LP_INDEX (_NDIS_ERROR_TYPEDEF_(0xC0350041L))
value ERROR_HV_INVALID_PARAMETER (_NDIS_ERROR_TYPEDEF_(0xC0350005L))
value ERROR_HV_INVALID_PARTITION_ID (_NDIS_ERROR_TYPEDEF_(0xC035000DL))
value ERROR_HV_INVALID_PARTITION_STATE (_NDIS_ERROR_TYPEDEF_(0xC0350007L))
value ERROR_HV_INVALID_PORT_ID (_NDIS_ERROR_TYPEDEF_(0xC0350011L))
value ERROR_HV_INVALID_PROXIMITY_DOMAIN_INFO (_NDIS_ERROR_TYPEDEF_(0xC035001AL))
value ERROR_HV_INVALID_REGISTER_VALUE (_NDIS_ERROR_TYPEDEF_(0xC0350050L))
value ERROR_HV_INVALID_SAVE_RESTORE_STATE (_NDIS_ERROR_TYPEDEF_(0xC0350017L))
value ERROR_HV_INVALID_SYNIC_STATE (_NDIS_ERROR_TYPEDEF_(0xC0350018L))
value ERROR_HV_INVALID_VP_INDEX (_NDIS_ERROR_TYPEDEF_(0xC035000EL))
value ERROR_HV_INVALID_VP_STATE (_NDIS_ERROR_TYPEDEF_(0xC0350015L))
value ERROR_HV_INVALID_VTL_STATE (_NDIS_ERROR_TYPEDEF_(0xC0350051L))
value ERROR_HV_MSR_ACCESS_FAILED (_NDIS_ERROR_TYPEDEF_(0xC0350080L))
value ERROR_HV_NESTED_VM_EXIT (_NDIS_ERROR_TYPEDEF_(0xC0350077L))
value ERROR_HV_NOT_ACKNOWLEDGED (_NDIS_ERROR_TYPEDEF_(0xC0350014L))
value ERROR_HV_NOT_ALLOWED_WITH_NESTED_VIRT_ACTIVE (_NDIS_ERROR_TYPEDEF_(0xC0350072L))
value ERROR_HV_NOT_PRESENT (_NDIS_ERROR_TYPEDEF_(0xC0351000L))
value ERROR_HV_NO_DATA (_NDIS_ERROR_TYPEDEF_(0xC035001BL))
value ERROR_HV_NO_RESOURCES (_NDIS_ERROR_TYPEDEF_(0xC035001DL))
value ERROR_HV_NX_NOT_DETECTED (_NDIS_ERROR_TYPEDEF_(0xC0350055L))
value ERROR_HV_OBJECT_IN_USE (_NDIS_ERROR_TYPEDEF_(0xC0350019L))
value ERROR_HV_OPERATION_DENIED (_NDIS_ERROR_TYPEDEF_(0xC0350008L))
value ERROR_HV_OPERATION_FAILED (_NDIS_ERROR_TYPEDEF_(0xC0350071L))
value ERROR_HV_PAGE_REQUEST_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0350060L))
value ERROR_HV_PARTITION_TOO_DEEP (_NDIS_ERROR_TYPEDEF_(0xC035000CL))
value ERROR_HV_PENDING_PAGE_REQUESTS (_NDIS_ERROR_TYPEDEF_(0x00350059L))
value ERROR_HV_PROCESSOR_STARTUP_TIMEOUT (_NDIS_ERROR_TYPEDEF_(0xC035003EL))
value ERROR_HV_PROPERTY_VALUE_OUT_OF_RANGE (_NDIS_ERROR_TYPEDEF_(0xC035000AL))
value ERROR_HV_SMX_ENABLED (_NDIS_ERROR_TYPEDEF_(0xC035003FL))
value ERROR_HV_UNKNOWN_PROPERTY (_NDIS_ERROR_TYPEDEF_(0xC0350009L))
value ERROR_HWNDS_HAVE_DIFF_PARENT (1441)
value ERROR_ICM_NOT_ENABLED (2018)
value ERROR_IEPORT_FULL (4341)
value ERROR_ILLEGAL_CHARACTER (582)
value ERROR_ILLEGAL_DLL_RELOCATION (623)
value ERROR_ILLEGAL_ELEMENT_ADDRESS (1162)
value ERROR_ILLEGAL_FLOAT_CONTEXT (579)
value ERROR_ILL_FORMED_PASSWORD (1324)
value ERROR_IMAGE_AT_DIFFERENT_BASE (807)
value ERROR_IMAGE_MACHINE_TYPE_MISMATCH (706)
value ERROR_IMAGE_MACHINE_TYPE_MISMATCH_EXE (720)
value ERROR_IMAGE_NOT_AT_BASE (700)
value ERROR_IMAGE_SUBSYSTEM_NOT_PRESENT (308)
value ERROR_IMPLEMENTATION_LIMIT (1292)
value ERROR_IMPLICIT_TRANSACTION_NOT_SUPPORTED (6725)
value ERROR_INCOMPATIBLE_SERVICE_PRIVILEGE (1297)
value ERROR_INCOMPATIBLE_SERVICE_SID_TYPE (1290)
value ERROR_INCOMPATIBLE_WITH_GLOBAL_SHORT_NAME_REGISTRY_SETTING (304)
value ERROR_INCORRECT_ACCOUNT_TYPE (8646)
value ERROR_INCORRECT_ADDRESS (1241)
value ERROR_INCORRECT_SIZE (1462)
value ERROR_INC_BACKUP (4003)
value ERROR_INDEX_ABSENT (1611)
value ERROR_INDEX_OUT_OF_BOUNDS (474)
value ERROR_INDIGENOUS_TYPE (4338)
value ERROR_INDOUBT_TRANSACTIONS_EXIST (6827)
value ERROR_INFLOOP_IN_RELOC_CHAIN (202)
value ERROR_INIT_STATUS_NEEDED (0x00000011)
value ERROR_INSTALL_ALREADY_RUNNING (1618)
value ERROR_INSTALL_CANCEL (15608)
value ERROR_INSTALL_DEREGISTRATION_FAILURE (15607)
value ERROR_INSTALL_FAILED (15609)
value ERROR_INSTALL_FAILURE (1603)
value ERROR_INSTALL_FIREWALL_SERVICE_NOT_RUNNING (15626)
value ERROR_INSTALL_FULLTRUST_HOSTRUNTIME_REQUIRES_MAIN_PACKAGE_FULLTRUST_CAPABILITY (15663)
value ERROR_INSTALL_INVALID_PACKAGE (15602)
value ERROR_INSTALL_INVALID_RELATED_SET_UPDATE (15639)
value ERROR_INSTALL_LANGUAGE_UNSUPPORTED (1623)
value ERROR_INSTALL_LOG_FAILURE (1622)
value ERROR_INSTALL_NETWORK_FAILURE (15605)
value ERROR_INSTALL_NOTUSED (1634)
value ERROR_INSTALL_OPEN_PACKAGE_FAILED (15600)
value ERROR_INSTALL_OPTIONAL_PACKAGE_APPLICATIONID_NOT_UNIQUE (15637)
value ERROR_INSTALL_OPTIONAL_PACKAGE_REQUIRES_MAIN_PACKAGE (15634)
value ERROR_INSTALL_OPTIONAL_PACKAGE_REQUIRES_MAIN_PACKAGE_FULLTRUST_CAPABILITY (15640)
value ERROR_INSTALL_OUT_OF_DISK_SPACE (15604)
value ERROR_INSTALL_PACKAGE_DOWNGRADE (15622)
value ERROR_INSTALL_PACKAGE_INVALID (1620)
value ERROR_INSTALL_PACKAGE_NOT_FOUND (15601)
value ERROR_INSTALL_PACKAGE_OPEN_FAILED (1619)
value ERROR_INSTALL_PACKAGE_REJECTED (1625)
value ERROR_INSTALL_PACKAGE_VERSION (1613)
value ERROR_INSTALL_PLATFORM_UNSUPPORTED (1633)
value ERROR_INSTALL_POLICY_FAILURE (15615)
value ERROR_INSTALL_PREREQUISITE_FAILED (15613)
value ERROR_INSTALL_REGISTRATION_FAILURE (15606)
value ERROR_INSTALL_REJECTED (1654)
value ERROR_INSTALL_REMOTE_DISALLOWED (1640)
value ERROR_INSTALL_REMOTE_PROHIBITED (1645)
value ERROR_INSTALL_RESOLVE_DEPENDENCY_FAILED (15603)
value ERROR_INSTALL_RESOLVE_HOSTRUNTIME_DEPENDENCY_FAILED (15665)
value ERROR_INSTALL_SERVICE_FAILURE (1601)
value ERROR_INSTALL_SERVICE_SAFEBOOT (1652)
value ERROR_INSTALL_SOURCE_ABSENT (1612)
value ERROR_INSTALL_SUSPEND (1604)
value ERROR_INSTALL_TEMP_UNWRITABLE (1632)
value ERROR_INSTALL_TRANSFORM_FAILURE (1624)
value ERROR_INSTALL_TRANSFORM_REJECTED (1644)
value ERROR_INSTALL_UI_FAILURE (1621)
value ERROR_INSTALL_USEREXIT (1602)
value ERROR_INSTALL_VOLUME_CORRUPT (15630)
value ERROR_INSTALL_VOLUME_NOT_EMPTY (15628)
value ERROR_INSTALL_VOLUME_OFFLINE (15629)
value ERROR_INSTALL_WRONG_PROCESSOR_ARCHITECTURE (15632)
value ERROR_INSTRUCTION_MISALIGNMENT (549)
value ERROR_INSUFFICIENT_BUFFER (122)
value ERROR_INSUFFICIENT_LOGON_INFO (608)
value ERROR_INSUFFICIENT_POWER (639)
value ERROR_INSUFFICIENT_RESOURCE_FOR_SPECIFIED_SHARED_SECTION_SIZE (781)
value ERROR_INSUFFICIENT_VIRTUAL_ADDR_RESOURCES (473)
value ERROR_INTERMIXED_KERNEL_EA_OPERATION (324)
value ERROR_INTERNAL_DB_CORRUPTION (1358)
value ERROR_INTERNAL_DB_ERROR (1383)
value ERROR_INTERNAL_ERROR (1359)
value ERROR_INTERRUPT_STILL_CONNECTED (764)
value ERROR_INTERRUPT_VECTOR_ALREADY_CONNECTED (763)
value ERROR_INVALID_ACCEL_HANDLE (1403)
value ERROR_INVALID_ACCESS (12)
value ERROR_INVALID_ACCOUNT_NAME (1315)
value ERROR_INVALID_ACE_CONDITION (805)
value ERROR_INVALID_ACL (1336)
value ERROR_INVALID_ADDRESS (487)
value ERROR_INVALID_AT_INTERRUPT_TIME (104)
value ERROR_INVALID_BLOCK (9)
value ERROR_INVALID_BLOCK_LENGTH (1106)
value ERROR_INVALID_CAP (320)
value ERROR_INVALID_CATEGORY (117)
value ERROR_INVALID_CLEANER (4310)
value ERROR_INVALID_CMM (2010)
value ERROR_INVALID_COLORINDEX (2022)
value ERROR_INVALID_COLORSPACE (2017)
value ERROR_INVALID_COMBOBOX_MESSAGE (1422)
value ERROR_INVALID_COMMAND_LINE (1639)
value ERROR_INVALID_COMPUTERNAME (1210)
value ERROR_INVALID_CRUNTIME_PARAMETER (1288)
value ERROR_INVALID_CURSOR_HANDLE (1402)
value ERROR_INVALID_DATA (13)
value ERROR_INVALID_DATATYPE (1804)
value ERROR_INVALID_DEVICE_OBJECT_PARAMETER (650)
value ERROR_INVALID_DLL (1154)
value ERROR_INVALID_DOMAINNAME (1212)
value ERROR_INVALID_DOMAIN_ROLE (1354)
value ERROR_INVALID_DOMAIN_STATE (1353)
value ERROR_INVALID_DRIVE (15)
value ERROR_INVALID_DRIVE_OBJECT (4321)
value ERROR_INVALID_DWP_HANDLE (1405)
value ERROR_INVALID_EA_HANDLE (278)
value ERROR_INVALID_EA_NAME (254)
value ERROR_INVALID_EDIT_HEIGHT (1424)
value ERROR_INVALID_ENVIRONMENT (1805)
value ERROR_INVALID_EVENTNAME (1211)
value ERROR_INVALID_EVENT_COUNT (151)
value ERROR_INVALID_EXCEPTION_HANDLER (310)
value ERROR_INVALID_EXE_SIGNATURE (191)
value ERROR_INVALID_FIELD (1616)
value ERROR_INVALID_FIELD_IN_PARAMETER_LIST (328)
value ERROR_INVALID_FILTER_PROC (1427)
value ERROR_INVALID_FLAGS (1004)
value ERROR_INVALID_FLAG_NUMBER (186)
value ERROR_INVALID_FORM_NAME (1902)
value ERROR_INVALID_FORM_SIZE (1903)
value ERROR_INVALID_FUNCTION (1)
value ERROR_INVALID_GROUPNAME (1209)
value ERROR_INVALID_GROUP_ATTRIBUTES (1345)
value ERROR_INVALID_GW_COMMAND (1443)
value ERROR_INVALID_HANDLE (6)
value ERROR_INVALID_HANDLE_STATE (1609)
value ERROR_INVALID_HOOK_FILTER (1426)
value ERROR_INVALID_HOOK_HANDLE (1404)
value ERROR_INVALID_HW_PROFILE (619)
value ERROR_INVALID_ICON_HANDLE (1414)
value ERROR_INVALID_ID_AUTHORITY (1343)
value ERROR_INVALID_IMAGE_HASH (577)
value ERROR_INVALID_IMPORT_OF_NON_DLL (1276)
value ERROR_INVALID_INDEX (1413)
value ERROR_INVALID_KERNEL_INFO_VERSION (340)
value ERROR_INVALID_KEYBOARD_HANDLE (1457)
value ERROR_INVALID_LABEL (1299)
value ERROR_INVALID_LB_MESSAGE (1432)
value ERROR_INVALID_LDT_DESCRIPTOR (564)
value ERROR_INVALID_LDT_OFFSET (563)
value ERROR_INVALID_LDT_SIZE (561)
value ERROR_INVALID_LEVEL (124)
value ERROR_INVALID_LIBRARY (4301)
value ERROR_INVALID_LIST_FORMAT (153)
value ERROR_INVALID_LOCK_RANGE (307)
value ERROR_INVALID_LOGON_HOURS (1328)
value ERROR_INVALID_LOGON_TYPE (1367)
value ERROR_INVALID_MEDIA (4300)
value ERROR_INVALID_MEDIA_POOL (4302)
value ERROR_INVALID_MEMBER (1388)
value ERROR_INVALID_MENU_HANDLE (1401)
value ERROR_INVALID_MESSAGE (1002)
value ERROR_INVALID_MESSAGEDEST (1218)
value ERROR_INVALID_MESSAGENAME (1217)
value ERROR_INVALID_MINALLOCSIZE (195)
value ERROR_INVALID_MODULETYPE (190)
value ERROR_INVALID_MONITOR_HANDLE (1461)
value ERROR_INVALID_MSGBOX_STYLE (1438)
value ERROR_INVALID_NAME (123)
value ERROR_INVALID_NETNAME (1214)
value ERROR_INVALID_OPERATION (4317)
value ERROR_INVALID_OPERATION_ON_QUORUM (5068)
value ERROR_INVALID_OPLOCK_PROTOCOL (301)
value ERROR_INVALID_ORDINAL (182)
value ERROR_INVALID_OWNER (1307)
value ERROR_INVALID_PACKAGE_SID_LENGTH (4253)
value ERROR_INVALID_PARAMETER (87)
value ERROR_INVALID_PASSWORD (86)
value ERROR_INVALID_PASSWORDNAME (1216)
value ERROR_INVALID_PATCH_XML (1650)
value ERROR_INVALID_PEP_INFO_VERSION (341)
value ERROR_INVALID_PIXEL_FORMAT (2000)
value ERROR_INVALID_PLUGPLAY_DEVICE_PATH (620)
value ERROR_INVALID_PORT_ATTRIBUTES (545)
value ERROR_INVALID_PRIMARY_GROUP (1308)
value ERROR_INVALID_PRINTER_COMMAND (1803)
value ERROR_INVALID_PRINTER_DRIVER_MANIFEST (3021)
value ERROR_INVALID_PRINTER_NAME (1801)
value ERROR_INVALID_PRINTER_STATE (1906)
value ERROR_INVALID_PRINT_MONITOR (3007)
value ERROR_INVALID_PRIORITY (1800)
value ERROR_INVALID_PROFILE (2011)
value ERROR_INVALID_QUOTA_LOWER (547)
value ERROR_INVALID_REPARSE_DATA (4392)
value ERROR_INVALID_RUNLEVEL_SETTING (15401)
value ERROR_INVALID_SCROLLBAR_RANGE (1448)
value ERROR_INVALID_SECURITY_DESCR (1338)
value ERROR_INVALID_SEGDPL (198)
value ERROR_INVALID_SEGMENT_NUMBER (180)
value ERROR_INVALID_SEPARATOR_FILE (1799)
value ERROR_INVALID_SERVER_STATE (1352)
value ERROR_INVALID_SERVICENAME (1213)
value ERROR_INVALID_SERVICE_ACCOUNT (1057)
value ERROR_INVALID_SERVICE_CONTROL (1052)
value ERROR_INVALID_SERVICE_LOCK (1071)
value ERROR_INVALID_SHARENAME (1215)
value ERROR_INVALID_SHOWWIN_COMMAND (1449)
value ERROR_INVALID_SID (1337)
value ERROR_INVALID_SIGNAL_NUMBER (209)
value ERROR_INVALID_SPI_VALUE (1439)
value ERROR_INVALID_STACKSEG (189)
value ERROR_INVALID_STAGED_SIGNATURE (15620)
value ERROR_INVALID_STARTING_CODESEG (188)
value ERROR_INVALID_STATE (5023)
value ERROR_INVALID_SUB_AUTHORITY (1335)
value ERROR_INVALID_TABLE (1628)
value ERROR_INVALID_TARGET_HANDLE (114)
value ERROR_INVALID_TASK_INDEX (1551)
value ERROR_INVALID_TASK_NAME (1550)
value ERROR_INVALID_THREAD_ID (1444)
value ERROR_INVALID_TIME (1901)
value ERROR_INVALID_TOKEN (315)
value ERROR_INVALID_TRANSACTION (6700)
value ERROR_INVALID_TRANSFORM (2020)
value ERROR_INVALID_UNWIND_TARGET (544)
value ERROR_INVALID_USER_BUFFER (1784)
value ERROR_INVALID_USER_PRINCIPAL_NAME (8636)
value ERROR_INVALID_VARIANT (604)
value ERROR_INVALID_VERIFY_SWITCH (118)
value ERROR_INVALID_WINDOW_HANDLE (1400)
value ERROR_INVALID_WINDOW_STYLE (2002)
value ERROR_INVALID_WORKSTATION (1329)
value ERROR_IOPL_NOT_ENABLED (197)
value ERROR_IO_DEVICE (1117)
value ERROR_IO_INCOMPLETE (996)
value ERROR_IO_PENDING (997)
value ERROR_IO_PREEMPTED (_HRESULT_TYPEDEF_(0x89010001L))
value ERROR_IO_PRIVILEGE_FAILED (571)
value ERROR_IO_REISSUE_AS_CACHED (3950)
value ERROR_IPSEC_AUTH_FIREWALL_DROP (13917)
value ERROR_IPSEC_BAD_SPI (13910)
value ERROR_IPSEC_CLEAR_TEXT_DROP (13916)
value ERROR_IPSEC_DEFAULT_MM_AUTH_NOT_FOUND (13014)
value ERROR_IPSEC_DEFAULT_MM_POLICY_NOT_FOUND (13013)
value ERROR_IPSEC_DEFAULT_QM_POLICY_NOT_FOUND (13015)
value ERROR_IPSEC_DOSP_BLOCK (13925)
value ERROR_IPSEC_DOSP_INVALID_PACKET (13927)
value ERROR_IPSEC_DOSP_KEYMOD_NOT_ALLOWED (13930)
value ERROR_IPSEC_DOSP_MAX_ENTRIES (13929)
value ERROR_IPSEC_DOSP_MAX_PER_IP_RATELIMIT_QUEUES (13932)
value ERROR_IPSEC_DOSP_NOT_INSTALLED (13931)
value ERROR_IPSEC_DOSP_RECEIVED_MULTICAST (13926)
value ERROR_IPSEC_DOSP_STATE_LOOKUP_FAILED (13928)
value ERROR_IPSEC_IKE_ADD_UPDATE_KEY_FAILED (13860)
value ERROR_IPSEC_IKE_ATTRIB_FAIL (13802)
value ERROR_IPSEC_IKE_AUTHORIZATION_FAILURE (13905)
value ERROR_IPSEC_IKE_AUTHORIZATION_FAILURE_WITH_OPTIONAL_RETRY (13907)
value ERROR_IPSEC_IKE_AUTH_FAIL (13801)
value ERROR_IPSEC_IKE_BENIGN_REINIT (13878)
value ERROR_IPSEC_IKE_CERT_CHAIN_POLICY_MISMATCH (13887)
value ERROR_IPSEC_IKE_CGA_AUTH_FAILED (13892)
value ERROR_IPSEC_IKE_COEXISTENCE_SUPPRESS (13902)
value ERROR_IPSEC_IKE_CRITICAL_PAYLOAD_NOT_RECOGNIZED (13823)
value ERROR_IPSEC_IKE_CRL_FAILED (13817)
value ERROR_IPSEC_IKE_DECRYPT (13867)
value ERROR_IPSEC_IKE_DH_FAIL (13822)
value ERROR_IPSEC_IKE_DH_FAILURE (13864)
value ERROR_IPSEC_IKE_DOS_COOKIE_SENT (13890)
value ERROR_IPSEC_IKE_DROP_NO_RESPONSE (13813)
value ERROR_IPSEC_IKE_ENCRYPT (13866)
value ERROR_IPSEC_IKE_ERROR (13816)
value ERROR_IPSEC_IKE_FAILQUERYSSP (13854)
value ERROR_IPSEC_IKE_FAILSSPINIT (13853)
value ERROR_IPSEC_IKE_GENERAL_PROCESSING_ERROR (13804)
value ERROR_IPSEC_IKE_GETSPIFAIL (13857)
value ERROR_IPSEC_IKE_INNER_IP_ASSIGNMENT_FAILURE (13899)
value ERROR_IPSEC_IKE_INVALID_AUTH_ALG (13874)
value ERROR_IPSEC_IKE_INVALID_AUTH_PAYLOAD (13889)
value ERROR_IPSEC_IKE_INVALID_CERT_KEYLEN (13881)
value ERROR_IPSEC_IKE_INVALID_CERT_TYPE (13819)
value ERROR_IPSEC_IKE_INVALID_COOKIE (13846)
value ERROR_IPSEC_IKE_INVALID_ENCRYPT_ALG (13873)
value ERROR_IPSEC_IKE_INVALID_FILTER (13858)
value ERROR_IPSEC_IKE_INVALID_GROUP (13865)
value ERROR_IPSEC_IKE_INVALID_HASH (13870)
value ERROR_IPSEC_IKE_INVALID_HASH_ALG (13871)
value ERROR_IPSEC_IKE_INVALID_HASH_SIZE (13872)
value ERROR_IPSEC_IKE_INVALID_HEADER (13824)
value ERROR_IPSEC_IKE_INVALID_KEY_USAGE (13818)
value ERROR_IPSEC_IKE_INVALID_MAJOR_VERSION (13880)
value ERROR_IPSEC_IKE_INVALID_MM_FOR_QM (13894)
value ERROR_IPSEC_IKE_INVALID_PAYLOAD (13843)
value ERROR_IPSEC_IKE_INVALID_POLICY (13861)
value ERROR_IPSEC_IKE_INVALID_RESPONDER_LIFETIME_NOTIFY (13879)
value ERROR_IPSEC_IKE_INVALID_SIG (13875)
value ERROR_IPSEC_IKE_INVALID_SIGNATURE (13826)
value ERROR_IPSEC_IKE_INVALID_SITUATION (13863)
value ERROR_IPSEC_IKE_KERBEROS_ERROR (13827)
value ERROR_IPSEC_IKE_KILL_DUMMY_NAP_TUNNEL (13898)
value ERROR_IPSEC_IKE_LOAD_FAILED (13876)
value ERROR_IPSEC_IKE_LOAD_SOFT_SA (13844)
value ERROR_IPSEC_IKE_MM_ACQUIRE_DROP (13809)
value ERROR_IPSEC_IKE_MM_DELAY_DROP (13814)
value ERROR_IPSEC_IKE_MM_EXPIRED (13885)
value ERROR_IPSEC_IKE_MM_LIMIT (13882)
value ERROR_IPSEC_IKE_NEGOTIATION_DISABLED (13883)
value ERROR_IPSEC_IKE_NEGOTIATION_PENDING (13803)
value ERROR_IPSEC_IKE_NEG_STATUS_BEGIN (13800)
value ERROR_IPSEC_IKE_NEG_STATUS_END (13897)
value ERROR_IPSEC_IKE_NEG_STATUS_EXTENDED_END (13909)
value ERROR_IPSEC_IKE_NOTCBPRIV (13851)
value ERROR_IPSEC_IKE_NO_CERT (13806)
value ERROR_IPSEC_IKE_NO_MM_POLICY (13850)
value ERROR_IPSEC_IKE_NO_PEER_CERT (13847)
value ERROR_IPSEC_IKE_NO_POLICY (13825)
value ERROR_IPSEC_IKE_NO_PRIVATE_KEY (13820)
value ERROR_IPSEC_IKE_NO_PUBLIC_KEY (13828)
value ERROR_IPSEC_IKE_OUT_OF_MEMORY (13859)
value ERROR_IPSEC_IKE_PEER_CRL_FAILED (13848)
value ERROR_IPSEC_IKE_PEER_DOESNT_SUPPORT_MOBIKE (13904)
value ERROR_IPSEC_IKE_PEER_MM_ASSUMED_INVALID (13886)
value ERROR_IPSEC_IKE_POLICY_CHANGE (13849)
value ERROR_IPSEC_IKE_POLICY_MATCH (13868)
value ERROR_IPSEC_IKE_PROCESS_ERR (13829)
value ERROR_IPSEC_IKE_PROCESS_ERR_CERT (13835)
value ERROR_IPSEC_IKE_PROCESS_ERR_CERT_REQ (13836)
value ERROR_IPSEC_IKE_PROCESS_ERR_DELETE (13841)
value ERROR_IPSEC_IKE_PROCESS_ERR_HASH (13837)
value ERROR_IPSEC_IKE_PROCESS_ERR_ID (13834)
value ERROR_IPSEC_IKE_PROCESS_ERR_KE (13833)
value ERROR_IPSEC_IKE_PROCESS_ERR_NATOA (13893)
value ERROR_IPSEC_IKE_PROCESS_ERR_NONCE (13839)
value ERROR_IPSEC_IKE_PROCESS_ERR_NOTIFY (13840)
value ERROR_IPSEC_IKE_PROCESS_ERR_PROP (13831)
value ERROR_IPSEC_IKE_PROCESS_ERR_SA (13830)
value ERROR_IPSEC_IKE_PROCESS_ERR_SIG (13838)
value ERROR_IPSEC_IKE_PROCESS_ERR_TRANS (13832)
value ERROR_IPSEC_IKE_PROCESS_ERR_VENDOR (13842)
value ERROR_IPSEC_IKE_QM_ACQUIRE_DROP (13810)
value ERROR_IPSEC_IKE_QM_DELAY_DROP (13815)
value ERROR_IPSEC_IKE_QM_EXPIRED (13895)
value ERROR_IPSEC_IKE_QM_LIMIT (13884)
value ERROR_IPSEC_IKE_QUEUE_DROP_MM (13811)
value ERROR_IPSEC_IKE_QUEUE_DROP_NO_MM (13812)
value ERROR_IPSEC_IKE_RATELIMIT_DROP (13903)
value ERROR_IPSEC_IKE_REQUIRE_CP_PAYLOAD_MISSING (13900)
value ERROR_IPSEC_IKE_RPC_DELETE (13877)
value ERROR_IPSEC_IKE_SA_DELETED (13807)
value ERROR_IPSEC_IKE_SA_REAPED (13808)
value ERROR_IPSEC_IKE_SECLOADFAIL (13852)
value ERROR_IPSEC_IKE_SHUTTING_DOWN (13891)
value ERROR_IPSEC_IKE_SIMULTANEOUS_REKEY (13821)
value ERROR_IPSEC_IKE_SOFT_SA_TORN_DOWN (13845)
value ERROR_IPSEC_IKE_SRVACQFAIL (13855)
value ERROR_IPSEC_IKE_SRVQUERYCRED (13856)
value ERROR_IPSEC_IKE_STRONG_CRED_AUTHORIZATION_AND_CERTMAP_FAILURE (13908)
value ERROR_IPSEC_IKE_STRONG_CRED_AUTHORIZATION_FAILURE (13906)
value ERROR_IPSEC_IKE_TIMED_OUT (13805)
value ERROR_IPSEC_IKE_TOO_MANY_FILTERS (13896)
value ERROR_IPSEC_IKE_UNEXPECTED_MESSAGE_ID (13888)
value ERROR_IPSEC_IKE_UNKNOWN_DOI (13862)
value ERROR_IPSEC_IKE_UNSUPPORTED_ID (13869)
value ERROR_IPSEC_INTEGRITY_CHECK_FAILED (13915)
value ERROR_IPSEC_INVALID_PACKET (13914)
value ERROR_IPSEC_KEY_MODULE_IMPERSONATION_NEGOTIATION_PENDING (13901)
value ERROR_IPSEC_MM_AUTH_EXISTS (13010)
value ERROR_IPSEC_MM_AUTH_IN_USE (13012)
value ERROR_IPSEC_MM_AUTH_NOT_FOUND (13011)
value ERROR_IPSEC_MM_AUTH_PENDING_DELETION (13022)
value ERROR_IPSEC_MM_FILTER_EXISTS (13006)
value ERROR_IPSEC_MM_FILTER_NOT_FOUND (13007)
value ERROR_IPSEC_MM_FILTER_PENDING_DELETION (13018)
value ERROR_IPSEC_MM_POLICY_EXISTS (13003)
value ERROR_IPSEC_MM_POLICY_IN_USE (13005)
value ERROR_IPSEC_MM_POLICY_NOT_FOUND (13004)
value ERROR_IPSEC_MM_POLICY_PENDING_DELETION (13021)
value ERROR_IPSEC_QM_POLICY_EXISTS (13000)
value ERROR_IPSEC_QM_POLICY_IN_USE (13002)
value ERROR_IPSEC_QM_POLICY_NOT_FOUND (13001)
value ERROR_IPSEC_QM_POLICY_PENDING_DELETION (13023)
value ERROR_IPSEC_REPLAY_CHECK_FAILED (13913)
value ERROR_IPSEC_SA_LIFETIME_EXPIRED (13911)
value ERROR_IPSEC_THROTTLE_DROP (13918)
value ERROR_IPSEC_TRANSPORT_FILTER_EXISTS (13008)
value ERROR_IPSEC_TRANSPORT_FILTER_NOT_FOUND (13009)
value ERROR_IPSEC_TRANSPORT_FILTER_PENDING_DELETION (13019)
value ERROR_IPSEC_TUNNEL_FILTER_EXISTS (13016)
value ERROR_IPSEC_TUNNEL_FILTER_NOT_FOUND (13017)
value ERROR_IPSEC_TUNNEL_FILTER_PENDING_DELETION (13020)
value ERROR_IPSEC_WRONG_SA (13912)
value ERROR_IRQ_BUSY (1119)
value ERROR_IS_JOINED (134)
value ERROR_IS_JOIN_PATH (147)
value ERROR_IS_JOIN_TARGET (133)
value ERROR_IS_SUBSTED (135)
value ERROR_IS_SUBST_PATH (146)
value ERROR_IS_SUBST_TARGET (149)
value ERROR_JOB_NO_CONTAINER (1505)
value ERROR_JOIN_TO_JOIN (138)
value ERROR_JOIN_TO_SUBST (140)
value ERROR_JOURNAL_DELETE_IN_PROGRESS (1178)
value ERROR_JOURNAL_ENTRY_DELETED (1181)
value ERROR_JOURNAL_HOOK_SET (1430)
value ERROR_JOURNAL_NOT_ACTIVE (1179)
value ERROR_KERNEL_APC (738)
value ERROR_KEY_DELETED (1018)
value ERROR_KEY_HAS_CHILDREN (1020)
value ERROR_KM_DRIVER_BLOCKED (1930)
value ERROR_LABEL_QUESTIONABLE (0x00000002)
value ERROR_LABEL_TOO_LONG (154)
value ERROR_LABEL_UNREADABLE (0x00000001)
value ERROR_LAST_ADMIN (1322)
value ERROR_LB_WITHOUT_TABSTOPS (1434)
value ERROR_LIBRARY_FULL (4322)
value ERROR_LIBRARY_OFFLINE (4305)
value ERROR_LICENSE_QUOTA_EXCEEDED (1395)
value ERROR_LINUX_SUBSYSTEM_NOT_PRESENT (414)
value ERROR_LINUX_SUBSYSTEM_UPDATE_REQUIRED (444)
value ERROR_LISTBOX_ID_NOT_FOUND (1416)
value ERROR_LM_CROSS_ENCRYPTION_REQUIRED (1390)
value ERROR_LOCAL_POLICY_MODIFICATION_NOT_SUPPORTED (8653)
value ERROR_LOCAL_USER_SESSION_KEY (1303)
value ERROR_LOCKED (212)
value ERROR_LOCK_FAILED (167)
value ERROR_LOCK_VIOLATION (33)
value ERROR_LOGIN_TIME_RESTRICTION (1239)
value ERROR_LOGIN_WKSTA_RESTRICTION (1240)
value ERROR_LOGON_FAILURE (1326)
value ERROR_LOGON_NOT_GRANTED (1380)
value ERROR_LOGON_SERVER_CONFLICT (568)
value ERROR_LOGON_SESSION_COLLISION (1366)
value ERROR_LOGON_SESSION_EXISTS (1363)
value ERROR_LOGON_TYPE_NOT_GRANTED (1385)
value ERROR_LOG_APPENDED_FLUSH_FAILED (6647)
value ERROR_LOG_ARCHIVE_IN_PROGRESS (6633)
value ERROR_LOG_ARCHIVE_NOT_IN_PROGRESS (6632)
value ERROR_LOG_BLOCKS_EXHAUSTED (6605)
value ERROR_LOG_BLOCK_INCOMPLETE (6603)
value ERROR_LOG_BLOCK_INVALID (6609)
value ERROR_LOG_BLOCK_VERSION (6608)
value ERROR_LOG_CANT_DELETE (6616)
value ERROR_LOG_CLIENT_ALREADY_REGISTERED (6636)
value ERROR_LOG_CLIENT_NOT_REGISTERED (6637)
value ERROR_LOG_CONTAINER_LIMIT_EXCEEDED (6617)
value ERROR_LOG_CONTAINER_OPEN_FAILED (6641)
value ERROR_LOG_CONTAINER_READ_FAILED (6639)
value ERROR_LOG_CONTAINER_STATE_INVALID (6642)
value ERROR_LOG_CONTAINER_WRITE_FAILED (6640)
value ERROR_LOG_CORRUPTION_DETECTED (6817)
value ERROR_LOG_DEDICATED (6631)
value ERROR_LOG_EPHEMERAL (6634)
value ERROR_LOG_FILE_FULL (1502)
value ERROR_LOG_FULL (6628)
value ERROR_LOG_FULL_HANDLER_IN_PROGRESS (6638)
value ERROR_LOG_GROWTH_FAILED (6833)
value ERROR_LOG_HARD_ERROR (718)
value ERROR_LOG_INCONSISTENT_SECURITY (6646)
value ERROR_LOG_INVALID_RANGE (6604)
value ERROR_LOG_METADATA_CORRUPT (6612)
value ERROR_LOG_METADATA_FLUSH_FAILED (6645)
value ERROR_LOG_METADATA_INCONSISTENT (6614)
value ERROR_LOG_METADATA_INVALID (6613)
value ERROR_LOG_MULTIPLEXED (6630)
value ERROR_LOG_NOT_ENOUGH_CONTAINERS (6635)
value ERROR_LOG_NO_RESTART (6611)
value ERROR_LOG_PINNED (6644)
value ERROR_LOG_PINNED_ARCHIVE_TAIL (6623)
value ERROR_LOG_PINNED_RESERVATION (6648)
value ERROR_LOG_POLICY_ALREADY_INSTALLED (6619)
value ERROR_LOG_POLICY_CONFLICT (6622)
value ERROR_LOG_POLICY_INVALID (6621)
value ERROR_LOG_POLICY_NOT_INSTALLED (6620)
value ERROR_LOG_READ_CONTEXT_INVALID (6606)
value ERROR_LOG_READ_MODE_INVALID (6610)
value ERROR_LOG_RECORDS_RESERVED_INVALID (6625)
value ERROR_LOG_RECORD_NONEXISTENT (6624)
value ERROR_LOG_RESERVATION_INVALID (6615)
value ERROR_LOG_RESIZE_INVALID_SIZE (6806)
value ERROR_LOG_RESTART_INVALID (6607)
value ERROR_LOG_SECTOR_INVALID (6600)
value ERROR_LOG_SECTOR_PARITY_INVALID (6601)
value ERROR_LOG_SECTOR_REMAPPED (6602)
value ERROR_LOG_SPACE_RESERVED_INVALID (6626)
value ERROR_LOG_START_OF_LOG (6618)
value ERROR_LOG_STATE_INVALID (6643)
value ERROR_LOG_TAIL_INVALID (6627)
value ERROR_LONGJUMP (682)
value ERROR_LOST_MODE_LOGON_RESTRICTION (1939)
value ERROR_LOST_WRITEBEHIND_DATA (596)
value ERROR_LOST_WRITEBEHIND_DATA_LOCAL_DISK_ERROR (790)
value ERROR_LOST_WRITEBEHIND_DATA_NETWORK_DISCONNECTED (788)
value ERROR_LOST_WRITEBEHIND_DATA_NETWORK_SERVER_ERROR (789)
value ERROR_LUIDS_EXHAUSTED (1334)
value ERROR_MACHINE_LOCKED (1271)
value ERROR_MACHINE_SCOPE_NOT_ALLOWED (15666)
value ERROR_MAGAZINE_NOT_PRESENT (1163)
value ERROR_MALFORMED_SUBSTITUTION_STRING (14094)
value ERROR_MAPPED_ALIGNMENT (1132)
value ERROR_MARKED_TO_DISALLOW_WRITES (348)
value ERROR_MARSHALL_OVERFLOW (603)
value ERROR_MAX_SESSIONS_REACHED (353)
value ERROR_MAX_THRDS_REACHED (164)
value ERROR_MCA_EXCEPTION (784)
value ERROR_MCA_INTERNAL_ERROR (15205)
value ERROR_MCA_INVALID_CAPABILITIES_STRING (15200)
value ERROR_MCA_INVALID_TECHNOLOGY_TYPE_RETURNED (15206)
value ERROR_MCA_INVALID_VCP_VERSION (15201)
value ERROR_MCA_MCCS_VERSION_MISMATCH (15203)
value ERROR_MCA_MONITOR_VIOLATES_MCCS_SPECIFICATION (15202)
value ERROR_MCA_OCCURED (651)
value ERROR_MCA_UNSUPPORTED_COLOR_TEMPERATURE (15207)
value ERROR_MCA_UNSUPPORTED_MCCS_VERSION (15204)
value ERROR_MEDIA_CHANGED (1110)
value ERROR_MEDIA_CHECK (679)
value ERROR_MEDIA_INCOMPATIBLE (4315)
value ERROR_MEDIA_NOT_AVAILABLE (4318)
value ERROR_MEDIA_OFFLINE (4304)
value ERROR_MEDIA_UNAVAILABLE (4308)
value ERROR_MEDIUM_NOT_ACCESSIBLE (4323)
value ERROR_MEMBERS_PRIMARY_GROUP (1374)
value ERROR_MEMBER_IN_ALIAS (1378)
value ERROR_MEMBER_IN_GROUP (1320)
value ERROR_MEMBER_NOT_IN_ALIAS (1377)
value ERROR_MEMBER_NOT_IN_GROUP (1321)
value ERROR_MEMORY_HARDWARE (779)
value ERROR_MENU_ITEM_NOT_FOUND (1456)
value ERROR_MESSAGE_EXCEEDS_MAX_SIZE (4336)
value ERROR_MESSAGE_SYNC_ONLY (1159)
value ERROR_METAFILE_NOT_SUPPORTED (2003)
value ERROR_META_EXPANSION_TOO_LONG (208)
value ERROR_MINIVERSION_INACCESSIBLE_FROM_SPECIFIED_TRANSACTION (6810)
value ERROR_MISSING_SYSTEMFILE (573)
value ERROR_MOD_NOT_FOUND (126)
value ERROR_MONITOR_INVALID_DESCRIPTOR_CHECKSUM (_HRESULT_TYPEDEF_(0xC0261003L))
value ERROR_MONITOR_INVALID_DETAILED_TIMING_BLOCK (_HRESULT_TYPEDEF_(0xC0261009L))
value ERROR_MONITOR_INVALID_MANUFACTURE_DATE (_HRESULT_TYPEDEF_(0xC026100AL))
value ERROR_MONITOR_INVALID_SERIAL_NUMBER_MONDSC_BLOCK (_HRESULT_TYPEDEF_(0xC0261006L))
value ERROR_MONITOR_INVALID_STANDARD_TIMING_BLOCK (_HRESULT_TYPEDEF_(0xC0261004L))
value ERROR_MONITOR_INVALID_USER_FRIENDLY_MONDSC_BLOCK (_HRESULT_TYPEDEF_(0xC0261007L))
value ERROR_MONITOR_NO_DESCRIPTOR (_HRESULT_TYPEDEF_(0x00261001L))
value ERROR_MONITOR_NO_MORE_DESCRIPTOR_DATA (_HRESULT_TYPEDEF_(0xC0261008L))
value ERROR_MONITOR_UNKNOWN_DESCRIPTOR_FORMAT (_HRESULT_TYPEDEF_(0x00261002L))
value ERROR_MONITOR_WMI_DATABLOCK_REGISTRATION_FAILED (_HRESULT_TYPEDEF_(0xC0261005L))
value ERROR_MORE_DATA (234)
value ERROR_MORE_WRITES (1120)
value ERROR_MOUNT_POINT_NOT_RESOLVED (649)
value ERROR_MP_PROCESSOR_MISMATCH (725)
value ERROR_MRM_AUTOMERGE_ENABLED (15139)
value ERROR_MRM_DIRECT_REF_TO_NON_DEFAULT_RESOURCE (15146)
value ERROR_MRM_DUPLICATE_ENTRY (15119)
value ERROR_MRM_DUPLICATE_MAP_NAME (15118)
value ERROR_MRM_FILEPATH_TOO_LONG (15121)
value ERROR_MRM_GENERATION_COUNT_MISMATCH (15147)
value ERROR_MRM_INDETERMINATE_QUALIFIER_VALUE (15138)
value ERROR_MRM_INVALID_FILE_TYPE (15112)
value ERROR_MRM_INVALID_PRICONFIG (15111)
value ERROR_MRM_INVALID_PRI_FILE (15126)
value ERROR_MRM_INVALID_QUALIFIER_OPERATOR (15137)
value ERROR_MRM_INVALID_QUALIFIER_VALUE (15114)
value ERROR_MRM_INVALID_RESOURCE_IDENTIFIER (15120)
value ERROR_MRM_MAP_NOT_FOUND (15135)
value ERROR_MRM_MISSING_DEFAULT_LANGUAGE (15160)
value ERROR_MRM_NAMED_RESOURCE_NOT_FOUND (15127)
value ERROR_MRM_NO_CANDIDATE (15115)
value ERROR_MRM_NO_CURRENT_VIEW_ON_THREAD (15143)
value ERROR_MRM_NO_MATCH_OR_DEFAULT_CANDIDATE (15116)
value ERROR_MRM_PACKAGE_NOT_FOUND (15159)
value ERROR_MRM_RESOURCE_TYPE_MISMATCH (15117)
value ERROR_MRM_RUNTIME_NO_DEFAULT_OR_NEUTRAL_RESOURCE (15110)
value ERROR_MRM_SCOPE_ITEM_CONFLICT (15161)
value ERROR_MRM_TOO_MANY_RESOURCES (15140)
value ERROR_MRM_UNKNOWN_QUALIFIER (15113)
value ERROR_MRM_UNSUPPORTED_DIRECTORY_TYPE (15122)
value ERROR_MRM_UNSUPPORTED_FILE_TYPE_FOR_LOAD_UNLOAD_PRI_FILE (15142)
value ERROR_MRM_UNSUPPORTED_FILE_TYPE_FOR_MERGE (15141)
value ERROR_MRM_UNSUPPORTED_PROFILE_TYPE (15136)
value ERROR_MR_MID_NOT_FOUND (317)
value ERROR_MUI_FILE_NOT_FOUND (15100)
value ERROR_MUI_FILE_NOT_LOADED (15105)
value ERROR_MUI_INTLSETTINGS_INVALID_LOCALE_NAME (15108)
value ERROR_MUI_INTLSETTINGS_UILANG_NOT_INSTALLED (15107)
value ERROR_MUI_INVALID_FILE (15101)
value ERROR_MUI_INVALID_LOCALE_NAME (15103)
value ERROR_MUI_INVALID_RC_CONFIG (15102)
value ERROR_MUI_INVALID_ULTIMATEFALLBACK_NAME (15104)
value ERROR_MULTIPLE_FAULT_VIOLATION (640)
value ERROR_MUTANT_LIMIT_EXCEEDED (587)
value ERROR_MUTUAL_AUTH_FAILED (1397)
value ERROR_NDIS_ADAPTER_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0x80340006L))
value ERROR_NDIS_ADAPTER_NOT_READY (_NDIS_ERROR_TYPEDEF_(0x80340011L))
value ERROR_NDIS_ADAPTER_REMOVED (_NDIS_ERROR_TYPEDEF_(0x80340018L))
value ERROR_NDIS_ALREADY_MAPPED (_NDIS_ERROR_TYPEDEF_(0x8034001DL))
value ERROR_NDIS_BAD_CHARACTERISTICS (_NDIS_ERROR_TYPEDEF_(0x80340005L))
value ERROR_NDIS_BAD_VERSION (_NDIS_ERROR_TYPEDEF_(0x80340004L))
value ERROR_NDIS_BUFFER_TOO_SHORT (_NDIS_ERROR_TYPEDEF_(0x80340016L))
value ERROR_NDIS_DEVICE_FAILED (_NDIS_ERROR_TYPEDEF_(0x80340008L))
value ERROR_NDIS_ERROR_READING_FILE (_NDIS_ERROR_TYPEDEF_(0x8034001CL))
value ERROR_NDIS_FILE_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0x8034001BL))
value ERROR_NDIS_GROUP_ADDRESS_IN_USE (_NDIS_ERROR_TYPEDEF_(0x8034001AL))
value ERROR_NDIS_INDICATION_REQUIRED (_NDIS_ERROR_TYPEDEF_(0x00340001L))
value ERROR_NDIS_INTERFACE_CLOSING (_NDIS_ERROR_TYPEDEF_(0x80340002L))
value ERROR_NDIS_INTERFACE_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0x8034002BL))
value ERROR_NDIS_INVALID_ADDRESS (_NDIS_ERROR_TYPEDEF_(0x80340022L))
value ERROR_NDIS_INVALID_DATA (_NDIS_ERROR_TYPEDEF_(0x80340015L))
value ERROR_NDIS_INVALID_DEVICE_REQUEST (_NDIS_ERROR_TYPEDEF_(0x80340010L))
value ERROR_NDIS_INVALID_LENGTH (_NDIS_ERROR_TYPEDEF_(0x80340014L))
value ERROR_NDIS_INVALID_OID (_NDIS_ERROR_TYPEDEF_(0x80340017L))
value ERROR_NDIS_INVALID_PACKET (_NDIS_ERROR_TYPEDEF_(0x8034000FL))
value ERROR_NDIS_INVALID_PORT (_NDIS_ERROR_TYPEDEF_(0x8034002DL))
value ERROR_NDIS_INVALID_PORT_STATE (_NDIS_ERROR_TYPEDEF_(0x8034002EL))
value ERROR_NDIS_LOW_POWER_STATE (_NDIS_ERROR_TYPEDEF_(0x8034002FL))
value ERROR_NDIS_MEDIA_DISCONNECTED (_NDIS_ERROR_TYPEDEF_(0x8034001FL))
value ERROR_NDIS_MULTICAST_EXISTS (_NDIS_ERROR_TYPEDEF_(0x8034000AL))
value ERROR_NDIS_MULTICAST_FULL (_NDIS_ERROR_TYPEDEF_(0x80340009L))
value ERROR_NDIS_MULTICAST_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0x8034000BL))
value ERROR_NDIS_NOT_SUPPORTED (_NDIS_ERROR_TYPEDEF_(0x803400BBL))
value ERROR_NDIS_NO_QUEUES (_NDIS_ERROR_TYPEDEF_(0x80340031L))
value ERROR_NDIS_OFFLOAD_CONNECTION_REJECTED (_NDIS_ERROR_TYPEDEF_(0xC0341012L))
value ERROR_NDIS_OFFLOAD_PATH_REJECTED (_NDIS_ERROR_TYPEDEF_(0xC0341013L))
value ERROR_NDIS_OFFLOAD_POLICY (_NDIS_ERROR_TYPEDEF_(0xC034100FL))
value ERROR_NDIS_OPEN_FAILED (_NDIS_ERROR_TYPEDEF_(0x80340007L))
value ERROR_NDIS_PAUSED (_NDIS_ERROR_TYPEDEF_(0x8034002AL))
value ERROR_NDIS_PM_PROTOCOL_OFFLOAD_LIST_FULL (_NDIS_ERROR_TYPEDEF_(0x80342004L))
value ERROR_NDIS_PM_WOL_PATTERN_LIST_FULL (_NDIS_ERROR_TYPEDEF_(0x80342003L))
value ERROR_NDIS_REINIT_REQUIRED (_NDIS_ERROR_TYPEDEF_(0x80340030L))
value ERROR_NDIS_REQUEST_ABORTED (_NDIS_ERROR_TYPEDEF_(0x8034000CL))
value ERROR_NDIS_RESET_IN_PROGRESS (_NDIS_ERROR_TYPEDEF_(0x8034000DL))
value ERROR_NDIS_RESOURCE_CONFLICT (_NDIS_ERROR_TYPEDEF_(0x8034001EL))
value ERROR_NDIS_UNSUPPORTED_MEDIA (_NDIS_ERROR_TYPEDEF_(0x80340019L))
value ERROR_NDIS_UNSUPPORTED_REVISION (_NDIS_ERROR_TYPEDEF_(0x8034002CL))
value ERROR_NEEDS_REGISTRATION (15631)
value ERROR_NEEDS_REMEDIATION (15612)
value ERROR_NEGATIVE_SEEK (131)
value ERROR_NESTING_NOT_ALLOWED (215)
value ERROR_NETLOGON_NOT_STARTED (1792)
value ERROR_NETNAME_DELETED (64)
value ERROR_NETWORK_ACCESS_DENIED (65)
value ERROR_NETWORK_ACCESS_DENIED_EDP (354)
value ERROR_NETWORK_AUTHENTICATION_PROMPT_CANCELED (3024)
value ERROR_NETWORK_BUSY (54)
value ERROR_NETWORK_NOT_AVAILABLE (5035)
value ERROR_NETWORK_UNREACHABLE (1231)
value ERROR_NET_OPEN_FAILED (570)
value ERROR_NET_WRITE_FAULT (88)
value ERROR_NOACCESS (998)
value ERROR_NODE_CANNOT_BE_CLUSTERED (5898)
value ERROR_NODE_CANT_HOST_RESOURCE (5071)
value ERROR_NODE_NOT_ACTIVE_CLUSTER_MEMBER (5980)
value ERROR_NODE_NOT_AVAILABLE (5036)
value ERROR_NOINTERFACE (632)
value ERROR_NOLOGON_INTERDOMAIN_TRUST_ACCOUNT (1807)
value ERROR_NOLOGON_SERVER_TRUST_ACCOUNT (1809)
value ERROR_NOLOGON_WORKSTATION_TRUST_ACCOUNT (1808)
value ERROR_NONCORE_GROUPS_FOUND (5937)
value ERROR_NONE_MAPPED (1332)
value ERROR_NONPAGED_SYSTEM_RESOURCES (1451)
value ERROR_NON_ACCOUNT_SID (1257)
value ERROR_NON_CSV_PATH (5950)
value ERROR_NON_DOMAIN_SID (1258)
value ERROR_NON_MDICHILD_WINDOW (1445)
value ERROR_NOTHING_TO_TERMINATE (758)
value ERROR_NOTIFICATION_GUID_ALREADY_DEFINED (309)
value ERROR_NOTIFY_CLEANUP (745)
value ERROR_NOTIFY_ENUM_DIR (1022)
value ERROR_NOT_ALLOWED_ON_SYSTEM_FILE (313)
value ERROR_NOT_ALL_ASSIGNED (1300)
value ERROR_NOT_APPCONTAINER (4250)
value ERROR_NOT_AUTHENTICATED (1244)
value ERROR_NOT_A_CLOUD_FILE (376)
value ERROR_NOT_A_CLOUD_SYNC_ROOT (405)
value ERROR_NOT_A_DAX_VOLUME (420)
value ERROR_NOT_A_REPARSE_POINT (4390)
value ERROR_NOT_A_TIERED_VOLUME (_HRESULT_TYPEDEF_(0x80830009L))
value ERROR_NOT_CAPABLE (775)
value ERROR_NOT_CHILD_WINDOW (1442)
value ERROR_NOT_CONNECTED (2250)
value ERROR_NOT_CONTAINER (1207)
value ERROR_NOT_DAX_MAPPABLE (421)
value ERROR_NOT_DOS_DISK (26)
value ERROR_NOT_EMPTY (4307)
value ERROR_NOT_ENOUGH_MEMORY (8)
value ERROR_NOT_ENOUGH_QUOTA (1816)
value ERROR_NOT_ENOUGH_SERVER_MEMORY (1130)
value ERROR_NOT_EXPORT_FORMAT (6008)
value ERROR_NOT_FOUND (1168)
value ERROR_NOT_GUI_PROCESS (1471)
value ERROR_NOT_JOINED (136)
value ERROR_NOT_LOCKED (158)
value ERROR_NOT_LOGGED_ON (1245)
value ERROR_NOT_LOGON_PROCESS (1362)
value ERROR_NOT_OWNER (288)
value ERROR_NOT_QUORUM_CAPABLE (5021)
value ERROR_NOT_QUORUM_CLASS (5025)
value ERROR_NOT_READY (21)
value ERROR_NOT_READ_FROM_COPY (337)
value ERROR_NOT_REDUNDANT_STORAGE (333)
value ERROR_NOT_REGISTRY_FILE (1017)
value ERROR_NOT_SAFEBOOT_SERVICE (1084)
value ERROR_NOT_SAFE_MODE_DRIVER (646)
value ERROR_NOT_SAME_DEVICE (17)
value ERROR_NOT_SAME_OBJECT (1656)
value ERROR_NOT_SNAPSHOT_VOLUME (6841)
value ERROR_NOT_SUBSTED (137)
value ERROR_NOT_SUPPORTED (50)
value ERROR_NOT_SUPPORTED_IN_APPCONTAINER (4252)
value ERROR_NOT_SUPPORTED_ON_DAX (360)
value ERROR_NOT_SUPPORTED_ON_SBS (1254)
value ERROR_NOT_SUPPORTED_ON_STANDARD_SERVER (8584)
value ERROR_NOT_SUPPORTED_WITH_AUDITING (499)
value ERROR_NOT_SUPPORTED_WITH_BTT (429)
value ERROR_NOT_SUPPORTED_WITH_BYPASSIO (493)
value ERROR_NOT_SUPPORTED_WITH_CACHED_HANDLE (509)
value ERROR_NOT_SUPPORTED_WITH_COMPRESSION (496)
value ERROR_NOT_SUPPORTED_WITH_DEDUPLICATION (498)
value ERROR_NOT_SUPPORTED_WITH_ENCRYPTION (495)
value ERROR_NOT_SUPPORTED_WITH_MONITORING (503)
value ERROR_NOT_SUPPORTED_WITH_REPLICATION (497)
value ERROR_NOT_SUPPORTED_WITH_SNAPSHOT (504)
value ERROR_NOT_SUPPORTED_WITH_VIRTUALIZATION (505)
value ERROR_NOT_TINY_STREAM (598)
value ERROR_NO_ACE_CONDITION (804)
value ERROR_NO_ADMIN_ACCESS_POINT (5090)
value ERROR_NO_APPLICABLE_APP_LICENSES_FOUND (_HRESULT_TYPEDEF_(0xC0EA0001L))
value ERROR_NO_ASSOCIATION (1155)
value ERROR_NO_BROWSER_SERVERS_FOUND (6118)
value ERROR_NO_BYPASSIO_DRIVER_SUPPORT (494)
value ERROR_NO_CALLBACK_ACTIVE (614)
value ERROR_NO_DATA (232)
value ERROR_NO_DATA_DETECTED (1104)
value ERROR_NO_EFS (6004)
value ERROR_NO_EVENT_PAIR (580)
value ERROR_NO_GUID_TRANSLATION (560)
value ERROR_NO_IMPERSONATION_TOKEN (1309)
value ERROR_NO_INHERITANCE (1391)
value ERROR_NO_LINK_TRACKING_IN_TRANSACTION (6852)
value ERROR_NO_LOGON_SERVERS (1311)
value ERROR_NO_LOG_SPACE (1019)
value ERROR_NO_MATCH (1169)
value ERROR_NO_MEDIA_IN_DRIVE (1112)
value ERROR_NO_MORE_DEVICES (1248)
value ERROR_NO_MORE_FILES (18)
value ERROR_NO_MORE_ITEMS (259)
value ERROR_NO_MORE_MATCHES (626)
value ERROR_NO_MORE_SEARCH_HANDLES (113)
value ERROR_NO_MORE_USER_HANDLES (1158)
value ERROR_NO_NETWORK (1222)
value ERROR_NO_NET_OR_BAD_PATH (1203)
value ERROR_NO_NVRAM_RESOURCES (1470)
value ERROR_NO_PAGEFILE (578)
value ERROR_NO_PHYSICALLY_ALIGNED_FREE_SPACE_FOUND (408)
value ERROR_NO_PROC_SLOTS (89)
value ERROR_NO_PROMOTION_ACTIVE (8222)
value ERROR_NO_QUOTAS_FOR_ACCOUNT (1302)
value ERROR_NO_RANGES_PROCESSED (312)
value ERROR_NO_RECOVERY_POLICY (6003)
value ERROR_NO_RECOVERY_PROGRAM (1082)
value ERROR_NO_SAVEPOINT_WITH_OPEN_FILES (6842)
value ERROR_NO_SCROLLBARS (1447)
value ERROR_NO_SECRETS (8620)
value ERROR_NO_SECURITY_ON_OBJECT (1350)
value ERROR_NO_SHUTDOWN_IN_PROGRESS (1116)
value ERROR_NO_SIGNAL_SENT (205)
value ERROR_NO_SITENAME (1919)
value ERROR_NO_SITE_SETTINGS_OBJECT (8619)
value ERROR_NO_SPOOL_SPACE (62)
value ERROR_NO_SUCH_ALIAS (1376)
value ERROR_NO_SUCH_DEVICE (433)
value ERROR_NO_SUCH_DOMAIN (1355)
value ERROR_NO_SUCH_GROUP (1319)
value ERROR_NO_SUCH_LOGON_SESSION (1312)
value ERROR_NO_SUCH_MEMBER (1387)
value ERROR_NO_SUCH_PACKAGE (1364)
value ERROR_NO_SUCH_PRIVILEGE (1313)
value ERROR_NO_SUCH_SITE (1249)
value ERROR_NO_SUCH_USER (1317)
value ERROR_NO_SUPPORTING_DRIVES (4339)
value ERROR_NO_SYSTEM_MENU (1437)
value ERROR_NO_SYSTEM_RESOURCES (1450)
value ERROR_NO_TASK_QUEUE (427)
value ERROR_NO_TOKEN (1008)
value ERROR_NO_TRACKING_SERVICE (1172)
value ERROR_NO_TRUST_LSA_SECRET (1786)
value ERROR_NO_TRUST_SAM_ACCOUNT (1787)
value ERROR_NO_TXF_METADATA (6816)
value ERROR_NO_UNICODE_TRANSLATION (1113)
value ERROR_NO_USER_KEYS (6006)
value ERROR_NO_USER_SESSION_KEY (1394)
value ERROR_NO_VOLUME_ID (1173)
value ERROR_NO_VOLUME_LABEL (125)
value ERROR_NO_WILDCARD_CHARACTERS (1417)
value ERROR_NO_WORK_DONE (235)
value ERROR_NO_WRITABLE_DC_FOUND (8621)
value ERROR_NO_YIELD_PERFORMED (721)
value ERROR_NTLM_BLOCKED (1937)
value ERROR_NT_CROSS_ENCRYPTION_REQUIRED (1386)
value ERROR_NULL_LM_PASSWORD (1304)
value ERROR_OBJECT_ALREADY_EXISTS (5010)
value ERROR_OBJECT_IN_LIST (5011)
value ERROR_OBJECT_IS_IMMUTABLE (4449)
value ERROR_OBJECT_NAME_EXISTS (698)
value ERROR_OBJECT_NOT_EXTERNALLY_BACKED (342)
value ERROR_OBJECT_NOT_FOUND (4312)
value ERROR_OBJECT_NO_LONGER_EXISTS (6807)
value ERROR_OFFLOAD_READ_FILE_NOT_SUPPORTED (4442)
value ERROR_OFFLOAD_READ_FLT_NOT_SUPPORTED (4440)
value ERROR_OFFLOAD_WRITE_FILE_NOT_SUPPORTED (4443)
value ERROR_OFFLOAD_WRITE_FLT_NOT_SUPPORTED (4441)
value ERROR_OFFSET_ALIGNMENT_VIOLATION (327)
value ERROR_OLD_WIN_VERSION (1150)
value ERROR_ONLY_IF_CONNECTED (1251)
value ERROR_OPEN_FAILED (110)
value ERROR_OPEN_FILES (2401)
value ERROR_OPERATION_ABORTED (995)
value ERROR_OPERATION_IN_PROGRESS (329)
value ERROR_OPERATION_NOT_ALLOWED_FROM_SYSTEM_COMPONENT (15145)
value ERROR_OPERATION_NOT_SUPPORTED_IN_TRANSACTION (6853)
value ERROR_OPLOCK_BREAK_IN_PROGRESS (742)
value ERROR_OPLOCK_HANDLE_CLOSED (803)
value ERROR_OPLOCK_NOT_GRANTED (300)
value ERROR_OPLOCK_SWITCHED_TO_NEW_HANDLE (800)
value ERROR_ORPHAN_NAME_EXHAUSTED (799)
value ERROR_OUTOFMEMORY (14)
value ERROR_OUT_OF_PAPER (28)
value ERROR_OUT_OF_STRUCTURES (84)
value ERROR_OVERRIDE_NOCHANGES (1252)
value ERROR_PACKAGED_SERVICE_REQUIRES_ADMIN_PRIVILEGES (15656)
value ERROR_PACKAGES_IN_USE (15618)
value ERROR_PACKAGES_REPUTATION_CHECK_FAILED (15643)
value ERROR_PACKAGES_REPUTATION_CHECK_TIMEDOUT (15644)
value ERROR_PACKAGE_ALREADY_EXISTS (15611)
value ERROR_PACKAGE_EXTERNAL_LOCATION_NOT_ALLOWED (15662)
value ERROR_PACKAGE_LACKS_CAPABILITY_FOR_MANDATORY_STARTUPTASKS (15664)
value ERROR_PACKAGE_LACKS_CAPABILITY_TO_DEPLOY_ON_HOST (15658)
value ERROR_PACKAGE_MOVE_BLOCKED_BY_STREAMING (15636)
value ERROR_PACKAGE_MOVE_FAILED (15627)
value ERROR_PACKAGE_NAME_MISMATCH (15670)
value ERROR_PACKAGE_NOT_REGISTERED_FOR_USER (15669)
value ERROR_PACKAGE_NOT_SUPPORTED_ON_FILESYSTEM (15635)
value ERROR_PACKAGE_REPOSITORY_CORRUPTED (15614)
value ERROR_PACKAGE_STAGING_ONHOLD (15638)
value ERROR_PACKAGE_UPDATING (15616)
value ERROR_PAGED_SYSTEM_RESOURCES (1452)
value ERROR_PAGEFILE_CREATE_FAILED (576)
value ERROR_PAGEFILE_NOT_SUPPORTED (491)
value ERROR_PAGEFILE_QUOTA (1454)
value ERROR_PAGEFILE_QUOTA_EXCEEDED (567)
value ERROR_PAGE_FAULT_COPY_ON_WRITE (749)
value ERROR_PAGE_FAULT_DEMAND_ZERO (748)
value ERROR_PAGE_FAULT_GUARD_PAGE (750)
value ERROR_PAGE_FAULT_PAGING_FILE (751)
value ERROR_PAGE_FAULT_TRANSITION (747)
value ERROR_PARAMETER_QUOTA_EXCEEDED (1283)
value ERROR_PARTIAL_COPY (299)
value ERROR_PARTITION_FAILURE (1105)
value ERROR_PARTITION_TERMINATING (1184)
value ERROR_PASSWORD_CHANGE_REQUIRED (1938)
value ERROR_PASSWORD_EXPIRED (1330)
value ERROR_PASSWORD_MUST_CHANGE (1907)
value ERROR_PASSWORD_RESTRICTION (1325)
value ERROR_PATCH_MANAGED_ADVERTISED_PRODUCT (1651)
value ERROR_PATCH_NO_SEQUENCE (1648)
value ERROR_PATCH_PACKAGE_INVALID (1636)
value ERROR_PATCH_PACKAGE_OPEN_FAILED (1635)
value ERROR_PATCH_PACKAGE_REJECTED (1643)
value ERROR_PATCH_PACKAGE_UNSUPPORTED (1637)
value ERROR_PATCH_REMOVAL_DISALLOWED (1649)
value ERROR_PATCH_REMOVAL_UNSUPPORTED (1646)
value ERROR_PATCH_TARGET_NOT_FOUND (1642)
value ERROR_PATH_BUSY (148)
value ERROR_PATH_NOT_FOUND (3)
value ERROR_PER_USER_TRUST_QUOTA_EXCEEDED (1932)
value ERROR_PIPE_BUSY (231)
value ERROR_PIPE_CONNECTED (535)
value ERROR_PIPE_LISTENING (536)
value ERROR_PIPE_LOCAL (229)
value ERROR_PIPE_NOT_CONNECTED (233)
value ERROR_PKINIT_FAILURE (1263)
value ERROR_PLATFORM_MANIFEST_BINARY_ID_NOT_FOUND (4574)
value ERROR_PLATFORM_MANIFEST_CATALOG_NOT_AUTHORIZED (4573)
value ERROR_PLATFORM_MANIFEST_FILE_NOT_AUTHORIZED (4572)
value ERROR_PLATFORM_MANIFEST_INVALID (4571)
value ERROR_PLATFORM_MANIFEST_NOT_ACTIVE (4575)
value ERROR_PLATFORM_MANIFEST_NOT_AUTHORIZED (4570)
value ERROR_PLATFORM_MANIFEST_NOT_SIGNED (4576)
value ERROR_PLUGPLAY_QUERY_VETOED (683)
value ERROR_PNP_BAD_MPS_TABLE (671)
value ERROR_PNP_INVALID_ID (674)
value ERROR_PNP_IRQ_TRANSLATION_FAILED (673)
value ERROR_PNP_QUERY_REMOVE_DEVICE_TIMEOUT (480)
value ERROR_PNP_QUERY_REMOVE_RELATED_DEVICE_TIMEOUT (481)
value ERROR_PNP_QUERY_REMOVE_UNRELATED_DEVICE_TIMEOUT (482)
value ERROR_PNP_REBOOT_REQUIRED (638)
value ERROR_PNP_RESTART_ENUMERATION (636)
value ERROR_PNP_TRANSLATION_FAILED (672)
value ERROR_POINT_NOT_FOUND (1171)
value ERROR_POLICY_OBJECT_NOT_FOUND (8219)
value ERROR_POLICY_ONLY_IN_DS (8220)
value ERROR_POPUP_ALREADY_ACTIVE (1446)
value ERROR_PORT_MESSAGE_TOO_LONG (546)
value ERROR_PORT_NOT_SET (642)
value ERROR_PORT_UNREACHABLE (1234)
value ERROR_POSSIBLE_DEADLOCK (1131)
value ERROR_POTENTIAL_FILE_FOUND (1180)
value ERROR_PREDEFINED_HANDLE (714)
value ERROR_PRIMARY_TRANSPORT_CONNECT_FAILED (746)
value ERROR_PRINTER_ALREADY_EXISTS (1802)
value ERROR_PRINTER_DELETED (1905)
value ERROR_PRINTER_DRIVER_ALREADY_INSTALLED (1795)
value ERROR_PRINTER_DRIVER_BLOCKED (3014)
value ERROR_PRINTER_DRIVER_DOWNLOAD_NEEDED (3019)
value ERROR_PRINTER_DRIVER_IN_USE (3001)
value ERROR_PRINTER_DRIVER_PACKAGE_IN_USE (3015)
value ERROR_PRINTER_DRIVER_WARNED (3013)
value ERROR_PRINTER_HAS_JOBS_QUEUED (3009)
value ERROR_PRINTER_NOT_FOUND (3012)
value ERROR_PRINTER_NOT_SHAREABLE (3022)
value ERROR_PRINTQ_FULL (61)
value ERROR_PRINT_CANCELLED (63)
value ERROR_PRINT_JOB_RESTART_REQUIRED (3020)
value ERROR_PRINT_MONITOR_ALREADY_INSTALLED (3006)
value ERROR_PRINT_MONITOR_IN_USE (3008)
value ERROR_PRINT_PROCESSOR_ALREADY_INSTALLED (3005)
value ERROR_PRIVATE_DIALOG_INDEX (1415)
value ERROR_PRIVILEGE_NOT_HELD (1314)
value ERROR_PRI_MERGE_ADD_FILE_FAILED (15151)
value ERROR_PRI_MERGE_BUNDLE_PACKAGES_NOT_ALLOWED (15155)
value ERROR_PRI_MERGE_INVALID_FILE_NAME (15158)
value ERROR_PRI_MERGE_LOAD_FILE_FAILED (15150)
value ERROR_PRI_MERGE_MAIN_PACKAGE_REQUIRED (15156)
value ERROR_PRI_MERGE_MISSING_SCHEMA (15149)
value ERROR_PRI_MERGE_MULTIPLE_MAIN_PACKAGES_NOT_ALLOWED (15154)
value ERROR_PRI_MERGE_MULTIPLE_PACKAGE_FAMILIES_NOT_ALLOWED (15153)
value ERROR_PRI_MERGE_RESOURCE_PACKAGE_REQUIRED (15157)
value ERROR_PRI_MERGE_VERSION_MISMATCH (15148)
value ERROR_PRI_MERGE_WRITE_FILE_FAILED (15152)
value ERROR_PROCESS_ABORTED (1067)
value ERROR_PROCESS_IN_JOB (760)
value ERROR_PROCESS_IS_PROTECTED (1293)
value ERROR_PROCESS_MODE_ALREADY_BACKGROUND (402)
value ERROR_PROCESS_MODE_NOT_BACKGROUND (403)
value ERROR_PROCESS_NOT_IN_JOB (759)
value ERROR_PROC_NOT_FOUND (127)
value ERROR_PRODUCT_UNINSTALLED (1614)
value ERROR_PRODUCT_VERSION (1638)
value ERROR_PROFILE_DOES_NOT_MATCH_DEVICE (2023)
value ERROR_PROFILE_NOT_ASSOCIATED_WITH_DEVICE (2015)
value ERROR_PROFILE_NOT_FOUND (2016)
value ERROR_PROFILING_AT_LIMIT (553)
value ERROR_PROFILING_NOT_STARTED (550)
value ERROR_PROFILING_NOT_STOPPED (551)
value ERROR_PROMOTION_ACTIVE (8221)
value ERROR_PROTOCOL_UNREACHABLE (1233)
value ERROR_PROVISION_OPTIONAL_PACKAGE_REQUIRES_MAIN_PACKAGE_PROVISIONED (15642)
value ERROR_PWD_HISTORY_CONFLICT (617)
value ERROR_PWD_TOO_LONG (657)
value ERROR_PWD_TOO_RECENT (616)
value ERROR_PWD_TOO_SHORT (615)
value ERROR_QUERY_STORAGE_ERROR (_NDIS_ERROR_TYPEDEF_(0x803A0001L))
value ERROR_QUIC_ALPN_NEG_FAILURE (_HRESULT_TYPEDEF_(0x80410007L))
value ERROR_QUIC_CONNECTION_IDLE (_HRESULT_TYPEDEF_(0x80410005L))
value ERROR_QUIC_CONNECTION_TIMEOUT (_HRESULT_TYPEDEF_(0x80410006L))
value ERROR_QUIC_HANDSHAKE_FAILURE (_HRESULT_TYPEDEF_(0x80410000L))
value ERROR_QUIC_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x80410003L))
value ERROR_QUIC_PROTOCOL_VIOLATION (_HRESULT_TYPEDEF_(0x80410004L))
value ERROR_QUIC_USER_CANCELED (_HRESULT_TYPEDEF_(0x80410002L))
value ERROR_QUIC_VER_NEG_FAILURE (_HRESULT_TYPEDEF_(0x80410001L))
value ERROR_QUORUMLOG_OPEN_FAILED (5028)
value ERROR_QUORUM_DISK_NOT_FOUND (5086)
value ERROR_QUORUM_NOT_ALLOWED_IN_THIS_GROUP (5928)
value ERROR_QUORUM_OWNER_ALIVE (5034)
value ERROR_QUORUM_RESOURCE (5020)
value ERROR_QUORUM_RESOURCE_ONLINE_FAILED (5027)
value ERROR_QUOTA_ACTIVITY (810)
value ERROR_QUOTA_LIST_INCONSISTENT (621)
value ERROR_RANGE_LIST_CONFLICT (627)
value ERROR_RANGE_NOT_FOUND (644)
value ERROR_RDP_PROTOCOL_ERROR (7065)
value ERROR_READ_FAULT (30)
value ERROR_RECEIVE_EXPEDITED (708)
value ERROR_RECEIVE_PARTIAL (707)
value ERROR_RECEIVE_PARTIAL_EXPEDITED (709)
value ERROR_RECOVERY_FAILURE (1279)
value ERROR_RECOVERY_FILE_CORRUPT (15619)
value ERROR_RECOVERY_NOT_NEEDED (6821)
value ERROR_REC_NON_EXISTENT (4005)
value ERROR_REDIRECTION_TO_DEFAULT_ACCOUNT_NOT_ALLOWED (15657)
value ERROR_REDIRECTOR_HAS_OPEN_HANDLES (1794)
value ERROR_REDIR_PAUSED (72)
value ERROR_REGISTRATION_FROM_REMOTE_DRIVE_NOT_SUPPORTED (15647)
value ERROR_REGISTRY_CORRUPT (1015)
value ERROR_REGISTRY_HIVE_RECOVERED (685)
value ERROR_REGISTRY_IO_FAILED (1016)
value ERROR_REGISTRY_QUOTA_LIMIT (613)
value ERROR_REGISTRY_RECOVERED (1014)
value ERROR_REG_NAT_CONSUMPTION (1261)
value ERROR_RELOC_CHAIN_XEEDS_SEGLIM (201)
value ERROR_REMOTE_FILE_VERSION_MISMATCH (6814)
value ERROR_REMOTE_PRINT_CONNECTIONS_BLOCKED (1936)
value ERROR_REMOTE_SESSION_LIMIT_EXCEEDED (1220)
value ERROR_REMOTE_STORAGE_MEDIA_ERROR (4352)
value ERROR_REMOTE_STORAGE_NOT_ACTIVE (4351)
value ERROR_REMOVE_FAILED (15610)
value ERROR_REM_NOT_LIST (51)
value ERROR_REPARSE (741)
value ERROR_REPARSE_ATTRIBUTE_CONFLICT (4391)
value ERROR_REPARSE_OBJECT (755)
value ERROR_REPARSE_POINT_ENCOUNTERED (4395)
value ERROR_REPARSE_TAG_INVALID (4393)
value ERROR_REPARSE_TAG_MISMATCH (4394)
value ERROR_REPLY_MESSAGE_MISMATCH (595)
value ERROR_REQUEST_ABORTED (1235)
value ERROR_REQUEST_OUT_OF_SEQUENCE (776)
value ERROR_REQUEST_PAUSED (3050)
value ERROR_REQUEST_REFUSED (4320)
value ERROR_REQUIRES_INTERACTIVE_WINDOWSTATION (1459)
value ERROR_REQ_NOT_ACCEP (71)
value ERROR_RESIDENT_FILE_NOT_SUPPORTED (334)
value ERROR_RESILIENCY_FILE_CORRUPT (15625)
value ERROR_RESMON_CREATE_FAILED (5017)
value ERROR_RESMON_INVALID_STATE (5084)
value ERROR_RESMON_ONLINE_FAILED (5018)
value ERROR_RESMON_SYSTEM_RESOURCES_LACKING (5956)
value ERROR_RESOURCEMANAGER_NOT_FOUND (6716)
value ERROR_RESOURCEMANAGER_READ_ONLY (6707)
value ERROR_RESOURCE_CALL_TIMED_OUT (5910)
value ERROR_RESOURCE_DATA_NOT_FOUND (1812)
value ERROR_RESOURCE_DISABLED (4309)
value ERROR_RESOURCE_ENUM_USER_STOP (15106)
value ERROR_RESOURCE_FAILED (5038)
value ERROR_RESOURCE_LANG_NOT_FOUND (1815)
value ERROR_RESOURCE_NAME_NOT_FOUND (1814)
value ERROR_RESOURCE_NOT_AVAILABLE (5006)
value ERROR_RESOURCE_NOT_FOUND (5007)
value ERROR_RESOURCE_NOT_IN_AVAILABLE_STORAGE (5965)
value ERROR_RESOURCE_NOT_ONLINE (5004)
value ERROR_RESOURCE_NOT_PRESENT (4316)
value ERROR_RESOURCE_ONLINE (5019)
value ERROR_RESOURCE_PROPERTIES_STORED (5024)
value ERROR_RESOURCE_PROPERTY_UNCHANGEABLE (5089)
value ERROR_RESOURCE_REQUIREMENTS_CHANGED (756)
value ERROR_RESOURCE_TYPE_NOT_FOUND (1813)
value ERROR_RESTART_APPLICATION (1467)
value ERROR_RESUME_HIBERNATION (727)
value ERROR_RETRY (1237)
value ERROR_RETURN_ADDRESS_HIJACK_ATTEMPT (1662)
value ERROR_REVISION_MISMATCH (1306)
value ERROR_RMODE_APP (1153)
value ERROR_RM_ALREADY_STARTED (6822)
value ERROR_RM_CANNOT_BE_FROZEN_FOR_SNAPSHOT (6728)
value ERROR_RM_DISCONNECTED (6819)
value ERROR_RM_METADATA_CORRUPT (6802)
value ERROR_RM_NOT_ACTIVE (6801)
value ERROR_ROLLBACK_TIMER_EXPIRED (6829)
value ERROR_ROWSNOTRELEASED (772)
value ERROR_RPL_NOT_ALLOWED (4006)
value ERROR_RUNLEVEL_SWITCH_AGENT_TIMEOUT (15403)
value ERROR_RUNLEVEL_SWITCH_IN_PROGRESS (15404)
value ERROR_RUNLEVEL_SWITCH_TIMEOUT (15402)
value ERROR_RWRAW_ENCRYPTED_FILE_NOT_ENCRYPTED (410)
value ERROR_RWRAW_ENCRYPTED_INVALID_EDATAINFO_FILEOFFSET (411)
value ERROR_RWRAW_ENCRYPTED_INVALID_EDATAINFO_FILERANGE (412)
value ERROR_RWRAW_ENCRYPTED_INVALID_EDATAINFO_PARAMETER (413)
value ERROR_RXACT_COMMITTED (744)
value ERROR_RXACT_COMMIT_FAILURE (1370)
value ERROR_RXACT_COMMIT_NECESSARY (678)
value ERROR_RXACT_INVALID_STATE (1369)
value ERROR_RXACT_STATE_CREATED (701)
value ERROR_SAME_DRIVE (143)
value ERROR_SAM_INIT_FAILURE (8541)
value ERROR_SCOPE_NOT_FOUND (318)
value ERROR_SCREEN_ALREADY_LOCKED (1440)
value ERROR_SCRUB_DATA_DISABLED (332)
value ERROR_SECCORE_INVALID_COMMAND (_HRESULT_TYPEDEF_(0xC0E80000L))
value ERROR_SECONDARY_IC_PROVIDER_NOT_REGISTERED (15321)
value ERROR_SECRET_TOO_LONG (1382)
value ERROR_SECTION_DIRECT_MAP_ONLY (819)
value ERROR_SECTOR_NOT_FOUND (27)
value ERROR_SECUREBOOT_FILE_REPLACED (4426)
value ERROR_SECUREBOOT_INVALID_POLICY (4422)
value ERROR_SECUREBOOT_NOT_BASE_POLICY (4434)
value ERROR_SECUREBOOT_NOT_ENABLED (4425)
value ERROR_SECUREBOOT_NOT_SUPPLEMENTAL_POLICY (4435)
value ERROR_SECUREBOOT_PLATFORM_ID_MISMATCH (4430)
value ERROR_SECUREBOOT_POLICY_MISSING_ANTIROLLBACKVERSION (4429)
value ERROR_SECUREBOOT_POLICY_NOT_AUTHORIZED (4427)
value ERROR_SECUREBOOT_POLICY_NOT_SIGNED (4424)
value ERROR_SECUREBOOT_POLICY_PUBLISHER_NOT_FOUND (4423)
value ERROR_SECUREBOOT_POLICY_ROLLBACK_DETECTED (4431)
value ERROR_SECUREBOOT_POLICY_UNKNOWN (4428)
value ERROR_SECUREBOOT_POLICY_UPGRADE_MISMATCH (4432)
value ERROR_SECUREBOOT_POLICY_VIOLATION (4421)
value ERROR_SECUREBOOT_REQUIRED_POLICY_FILE_MISSING (4433)
value ERROR_SECUREBOOT_ROLLBACK_DETECTED (4420)
value ERROR_SECURITY_DENIES_OPERATION (447)
value ERROR_SECURITY_STREAM_IS_INCONSISTENT (306)
value ERROR_SEEK (25)
value ERROR_SEEK_ON_DEVICE (132)
value ERROR_SEGMENT_NOTIFICATION (702)
value ERROR_SEM_IS_SET (102)
value ERROR_SEM_NOT_FOUND (187)
value ERROR_SEM_OWNER_DIED (105)
value ERROR_SEM_TIMEOUT (121)
value ERROR_SEM_USER_LIMIT (106)
value ERROR_SERIAL_NO_DEVICE (1118)
value ERROR_SERVER_DISABLED (1341)
value ERROR_SERVER_HAS_OPEN_HANDLES (1811)
value ERROR_SERVER_NOT_DISABLED (1342)
value ERROR_SERVER_SHUTDOWN_IN_PROGRESS (1255)
value ERROR_SERVER_SID_MISMATCH (628)
value ERROR_SERVER_TRANSPORT_CONFLICT (816)
value ERROR_SERVICES_FAILED_AUTOSTART (15405)
value ERROR_SERVICE_ALREADY_RUNNING (1056)
value ERROR_SERVICE_CANNOT_ACCEPT_CTRL (1061)
value ERROR_SERVICE_DATABASE_LOCKED (1055)
value ERROR_SERVICE_DEPENDENCY_DELETED (1075)
value ERROR_SERVICE_DEPENDENCY_FAIL (1068)
value ERROR_SERVICE_DISABLED (1058)
value ERROR_SERVICE_DOES_NOT_EXIST (1060)
value ERROR_SERVICE_EXISTS (1073)
value ERROR_SERVICE_EXISTS_AS_NON_PACKAGED_SERVICE (15655)
value ERROR_SERVICE_LOGON_FAILED (1069)
value ERROR_SERVICE_MARKED_FOR_DELETE (1072)
value ERROR_SERVICE_NEVER_STARTED (1077)
value ERROR_SERVICE_NOTIFICATION (716)
value ERROR_SERVICE_NOTIFY_CLIENT_LAGGING (1294)
value ERROR_SERVICE_NOT_ACTIVE (1062)
value ERROR_SERVICE_NOT_FOUND (1243)
value ERROR_SERVICE_NOT_IN_EXE (1083)
value ERROR_SERVICE_NO_THREAD (1054)
value ERROR_SERVICE_REQUEST_TIMEOUT (1053)
value ERROR_SERVICE_SPECIFIC_ERROR (1066)
value ERROR_SERVICE_START_HANG (1070)
value ERROR_SESSION_CREDENTIAL_CONFLICT (1219)
value ERROR_SESSION_KEY_TOO_SHORT (501)
value ERROR_SETCOUNT_ON_BAD_LB (1433)
value ERROR_SETMARK_DETECTED (1103)
value ERROR_SET_CONTEXT_DENIED (1660)
value ERROR_SET_NOT_FOUND (1170)
value ERROR_SET_POWER_STATE_FAILED (1141)
value ERROR_SET_POWER_STATE_VETOED (1140)
value ERROR_SEVERITY_ERROR (0xC0000000)
value ERROR_SEVERITY_INFORMATIONAL (0x40000000)
value ERROR_SEVERITY_SUCCESS (0x00000000)
value ERROR_SEVERITY_WARNING (0x80000000)
value ERROR_SHARED_POLICY (8218)
value ERROR_SHARING_BUFFER_EXCEEDED (36)
value ERROR_SHARING_PAUSED (70)
value ERROR_SHARING_VIOLATION (32)
value ERROR_SHORT_NAMES_NOT_ENABLED_ON_VOLUME (305)
value ERROR_SHUTDOWN_CLUSTER (5008)
value ERROR_SHUTDOWN_DISKS_NOT_IN_MAINTENANCE_MODE (1192)
value ERROR_SHUTDOWN_IN_PROGRESS (1115)
value ERROR_SHUTDOWN_IS_SCHEDULED (1190)
value ERROR_SHUTDOWN_USERS_LOGGED_ON (1191)
value ERROR_SIGNAL_PENDING (162)
value ERROR_SIGNAL_REFUSED (156)
value ERROR_SIGNED_PACKAGE_INVALID_PUBLISHER_NAMESPACE (15661)
value ERROR_SINGLETON_RESOURCE_INSTALLED_IN_ACTIVE_USER (15653)
value ERROR_SINGLE_INSTANCE_APP (1152)
value ERROR_SLOT_NOT_PRESENT (0x00000004)
value ERROR_SMARTCARD_SUBSYSTEM_FAILURE (1264)
value ERROR_SMB_BAD_CLUSTER_DIALECT (_HRESULT_TYPEDEF_(0xC05D0001L))
value ERROR_SMB_GUEST_LOGON_BLOCKED (1272)
value ERROR_SMB_NO_PREAUTH_INTEGRITY_HASH_OVERLAP (_HRESULT_TYPEDEF_(0xC05D0000L))
value ERROR_SMB_NO_SIGNING_ALGORITHM_OVERLAP (_HRESULT_TYPEDEF_(0xC05D0002L))
value ERROR_SMI_PRIMITIVE_INSTALLER_FAILED (14108)
value ERROR_SMR_GARBAGE_COLLECTION_REQUIRED (4445)
value ERROR_SOME_NOT_MAPPED (1301)
value ERROR_SOURCE_ELEMENT_EMPTY (1160)
value ERROR_SPACES_ALLOCATION_SIZE_INVALID (_HRESULT_TYPEDEF_(0x80E7000EL))
value ERROR_SPACES_CACHE_FULL (_HRESULT_TYPEDEF_(0x80E70026L))
value ERROR_SPACES_CORRUPT_METADATA (_HRESULT_TYPEDEF_(0x80E70018L))
value ERROR_SPACES_DRIVE_LOST_DATA (_HRESULT_TYPEDEF_(0x80E7001FL))
value ERROR_SPACES_DRIVE_NOT_READY (_HRESULT_TYPEDEF_(0x80E7001DL))
value ERROR_SPACES_DRIVE_OPERATIONAL_STATE_INVALID (_HRESULT_TYPEDEF_(0x80E70012L))
value ERROR_SPACES_DRIVE_REDUNDANCY_INVALID (_HRESULT_TYPEDEF_(0x80E70006L))
value ERROR_SPACES_DRIVE_SECTOR_SIZE_INVALID (_HRESULT_TYPEDEF_(0x80E70004L))
value ERROR_SPACES_DRIVE_SPLIT (_HRESULT_TYPEDEF_(0x80E7001EL))
value ERROR_SPACES_DRT_FULL (_HRESULT_TYPEDEF_(0x80E70019L))
value ERROR_SPACES_ENCLOSURE_AWARE_INVALID (_HRESULT_TYPEDEF_(0x80E7000FL))
value ERROR_SPACES_ENTRY_INCOMPLETE (_HRESULT_TYPEDEF_(0x80E70013L))
value ERROR_SPACES_ENTRY_INVALID (_HRESULT_TYPEDEF_(0x80E70014L))
value ERROR_SPACES_EXTENDED_ERROR (_HRESULT_TYPEDEF_(0x80E7000CL))
value ERROR_SPACES_FAULT_DOMAIN_TYPE_INVALID (_HRESULT_TYPEDEF_(0x80E70001L))
value ERROR_SPACES_FLUSH_METADATA (_HRESULT_TYPEDEF_(0x80E70025L))
value ERROR_SPACES_INCONSISTENCY (_HRESULT_TYPEDEF_(0x80E7001AL))
value ERROR_SPACES_INTERLEAVE_LENGTH_INVALID (_HRESULT_TYPEDEF_(0x80E70009L))
value ERROR_SPACES_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x80E70002L))
value ERROR_SPACES_LOG_NOT_READY (_HRESULT_TYPEDEF_(0x80E7001BL))
value ERROR_SPACES_MAP_REQUIRED (_HRESULT_TYPEDEF_(0x80E70016L))
value ERROR_SPACES_MARK_DIRTY (_HRESULT_TYPEDEF_(0x80E70020L))
value ERROR_SPACES_NOT_ENOUGH_DRIVES (_HRESULT_TYPEDEF_(0x80E7000BL))
value ERROR_SPACES_NO_REDUNDANCY (_HRESULT_TYPEDEF_(0x80E7001CL))
value ERROR_SPACES_NUMBER_OF_COLUMNS_INVALID (_HRESULT_TYPEDEF_(0x80E7000AL))
value ERROR_SPACES_NUMBER_OF_DATA_COPIES_INVALID (_HRESULT_TYPEDEF_(0x80E70007L))
value ERROR_SPACES_NUMBER_OF_GROUPS_INVALID (_HRESULT_TYPEDEF_(0x80E70011L))
value ERROR_SPACES_PARITY_LAYOUT_INVALID (_HRESULT_TYPEDEF_(0x80E70008L))
value ERROR_SPACES_POOL_WAS_DELETED (_HRESULT_TYPEDEF_(0x00E70001L))
value ERROR_SPACES_PROVISIONING_TYPE_INVALID (_HRESULT_TYPEDEF_(0x80E7000DL))
value ERROR_SPACES_REPAIR_IN_PROGRESS (_HRESULT_TYPEDEF_(0x80E70027L))
value ERROR_SPACES_RESILIENCY_TYPE_INVALID (_HRESULT_TYPEDEF_(0x80E70003L))
value ERROR_SPACES_UNSUPPORTED_VERSION (_HRESULT_TYPEDEF_(0x80E70017L))
value ERROR_SPACES_UPDATE_COLUMN_STATE (_HRESULT_TYPEDEF_(0x80E70015L))
value ERROR_SPACES_WRITE_CACHE_SIZE_INVALID (_HRESULT_TYPEDEF_(0x80E70010L))
value ERROR_SPARSE_FILE_NOT_SUPPORTED (490)
value ERROR_SPARSE_NOT_ALLOWED_IN_TRANSACTION (6844)
value ERROR_SPECIAL_ACCOUNT (1371)
value ERROR_SPECIAL_GROUP (1372)
value ERROR_SPECIAL_USER (1373)
value ERROR_SPL_NO_ADDJOB (3004)
value ERROR_SPL_NO_STARTDOC (3003)
value ERROR_SPOOL_FILE_NOT_FOUND (3002)
value ERROR_SRC_SRV_DLL_LOAD_FAILED (428)
value ERROR_STACK_BUFFER_OVERRUN (1282)
value ERROR_STACK_OVERFLOW (1001)
value ERROR_STACK_OVERFLOW_READ (599)
value ERROR_STAGEFROMUPDATEAGENT_PACKAGE_NOT_APPLICABLE (15668)
value ERROR_STATE_COMPOSITE_SETTING_VALUE_SIZE_LIMIT_EXCEEDED (15815)
value ERROR_STATE_CONTAINER_NAME_SIZE_LIMIT_EXCEEDED (15818)
value ERROR_STATE_CREATE_CONTAINER_FAILED (15805)
value ERROR_STATE_DELETE_CONTAINER_FAILED (15806)
value ERROR_STATE_DELETE_SETTING_FAILED (15809)
value ERROR_STATE_ENUMERATE_CONTAINER_FAILED (15813)
value ERROR_STATE_ENUMERATE_SETTINGS_FAILED (15814)
value ERROR_STATE_GET_VERSION_FAILED (15801)
value ERROR_STATE_LOAD_STORE_FAILED (15800)
value ERROR_STATE_OPEN_CONTAINER_FAILED (15804)
value ERROR_STATE_QUERY_SETTING_FAILED (15810)
value ERROR_STATE_READ_COMPOSITE_SETTING_FAILED (15811)
value ERROR_STATE_READ_SETTING_FAILED (15807)
value ERROR_STATE_SETTING_NAME_SIZE_LIMIT_EXCEEDED (15817)
value ERROR_STATE_SETTING_VALUE_SIZE_LIMIT_EXCEEDED (15816)
value ERROR_STATE_SET_VERSION_FAILED (15802)
value ERROR_STATE_STRUCTURED_RESET_FAILED (15803)
value ERROR_STATE_WRITE_COMPOSITE_SETTING_FAILED (15812)
value ERROR_STATE_WRITE_SETTING_FAILED (15808)
value ERROR_STATIC_INIT (4002)
value ERROR_STOPPED_ON_SYMLINK (681)
value ERROR_STORAGE_LOST_DATA_PERSISTENCE (368)
value ERROR_STORAGE_RESERVE_ALREADY_EXISTS (418)
value ERROR_STORAGE_RESERVE_DOES_NOT_EXIST (417)
value ERROR_STORAGE_RESERVE_ID_INVALID (416)
value ERROR_STORAGE_RESERVE_NOT_EMPTY (419)
value ERROR_STORAGE_STACK_ACCESS_DENIED (472)
value ERROR_STORAGE_TOPOLOGY_ID_MISMATCH (345)
value ERROR_STREAM_MINIVERSION_NOT_FOUND (6808)
value ERROR_STREAM_MINIVERSION_NOT_VALID (6809)
value ERROR_STRICT_CFG_VIOLATION (1657)
value ERROR_SUBST_TO_JOIN (141)
value ERROR_SUBST_TO_SUBST (139)
value ERROR_SUCCESS (0)
value ERROR_SUCCESS_REBOOT_INITIATED (1641)
value ERROR_SUCCESS_REBOOT_REQUIRED (3010)
value ERROR_SUCCESS_RESTART_REQUIRED (3011)
value ERROR_SVHDX_ERROR_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0xC05CFF00L))
value ERROR_SVHDX_ERROR_STORED (_HRESULT_TYPEDEF_(0xC05C0000L))
value ERROR_SVHDX_NO_INITIATOR (_HRESULT_TYPEDEF_(0xC05CFF0BL))
value ERROR_SVHDX_RESERVATION_CONFLICT (_HRESULT_TYPEDEF_(0xC05CFF07L))
value ERROR_SVHDX_UNIT_ATTENTION_AVAILABLE (_HRESULT_TYPEDEF_(0xC05CFF01L))
value ERROR_SVHDX_UNIT_ATTENTION_CAPACITY_DATA_CHANGED (_HRESULT_TYPEDEF_(0xC05CFF02L))
value ERROR_SVHDX_UNIT_ATTENTION_OPERATING_DEFINITION_CHANGED (_HRESULT_TYPEDEF_(0xC05CFF06L))
value ERROR_SVHDX_UNIT_ATTENTION_REGISTRATIONS_PREEMPTED (_HRESULT_TYPEDEF_(0xC05CFF05L))
value ERROR_SVHDX_UNIT_ATTENTION_RESERVATIONS_PREEMPTED (_HRESULT_TYPEDEF_(0xC05CFF03L))
value ERROR_SVHDX_UNIT_ATTENTION_RESERVATIONS_RELEASED (_HRESULT_TYPEDEF_(0xC05CFF04L))
value ERROR_SVHDX_VERSION_MISMATCH (_HRESULT_TYPEDEF_(0xC05CFF09L))
value ERROR_SVHDX_WRONG_FILE_TYPE (_HRESULT_TYPEDEF_(0xC05CFF08L))
value ERROR_SWAPERROR (999)
value ERROR_SXS_ACTIVATION_CONTEXT_DISABLED (14006)
value ERROR_SXS_ASSEMBLY_IS_NOT_A_DEPLOYMENT (14103)
value ERROR_SXS_ASSEMBLY_MISSING (14081)
value ERROR_SXS_ASSEMBLY_NOT_FOUND (14003)
value ERROR_SXS_ASSEMBLY_NOT_LOCKED (14097)
value ERROR_SXS_CANT_GEN_ACTCTX (14001)
value ERROR_SXS_COMPONENT_STORE_CORRUPT (14098)
value ERROR_SXS_CORRUPTION (14083)
value ERROR_SXS_CORRUPT_ACTIVATION_STACK (14082)
value ERROR_SXS_DUPLICATE_ACTIVATABLE_CLASS (14111)
value ERROR_SXS_DUPLICATE_ASSEMBLY_NAME (14027)
value ERROR_SXS_DUPLICATE_CLSID (14023)
value ERROR_SXS_DUPLICATE_DLL_NAME (14021)
value ERROR_SXS_DUPLICATE_IID (14024)
value ERROR_SXS_DUPLICATE_PROGID (14026)
value ERROR_SXS_DUPLICATE_TLBID (14025)
value ERROR_SXS_DUPLICATE_WINDOWCLASS_NAME (14022)
value ERROR_SXS_EARLY_DEACTIVATION (14084)
value ERROR_SXS_FILE_HASH_MISMATCH (14028)
value ERROR_SXS_FILE_HASH_MISSING (14110)
value ERROR_SXS_FILE_NOT_PART_OF_ASSEMBLY (14104)
value ERROR_SXS_IDENTITIES_DIFFERENT (14102)
value ERROR_SXS_IDENTITY_DUPLICATE_ATTRIBUTE (14092)
value ERROR_SXS_IDENTITY_PARSE_ERROR (14093)
value ERROR_SXS_INCORRECT_PUBLIC_KEY_TOKEN (14095)
value ERROR_SXS_INVALID_ACTCTXDATA_FORMAT (14002)
value ERROR_SXS_INVALID_ASSEMBLY_IDENTITY_ATTRIBUTE (14017)
value ERROR_SXS_INVALID_ASSEMBLY_IDENTITY_ATTRIBUTE_NAME (14080)
value ERROR_SXS_INVALID_DEACTIVATION (14085)
value ERROR_SXS_INVALID_IDENTITY_ATTRIBUTE_NAME (14091)
value ERROR_SXS_INVALID_IDENTITY_ATTRIBUTE_VALUE (14090)
value ERROR_SXS_INVALID_XML_NAMESPACE_URI (14014)
value ERROR_SXS_KEY_NOT_FOUND (14007)
value ERROR_SXS_LEAF_MANIFEST_DEPENDENCY_NOT_INSTALLED (14016)
value ERROR_SXS_MANIFEST_FORMAT_ERROR (14004)
value ERROR_SXS_MANIFEST_IDENTITY_SAME_BUT_CONTENTS_DIFFERENT (14101)
value ERROR_SXS_MANIFEST_INVALID_REQUIRED_DEFAULT_NAMESPACE (14019)
value ERROR_SXS_MANIFEST_MISSING_REQUIRED_DEFAULT_NAMESPACE (14018)
value ERROR_SXS_MANIFEST_PARSE_ERROR (14005)
value ERROR_SXS_MANIFEST_TOO_BIG (14105)
value ERROR_SXS_MISSING_ASSEMBLY_IDENTITY_ATTRIBUTE (14079)
value ERROR_SXS_MULTIPLE_DEACTIVATION (14086)
value ERROR_SXS_POLICY_PARSE_ERROR (14029)
value ERROR_SXS_PRIVATE_MANIFEST_CROSS_PATH_WITH_REPARSE_POINT (14020)
value ERROR_SXS_PROCESS_DEFAULT_ALREADY_SET (14011)
value ERROR_SXS_PROCESS_TERMINATION_REQUESTED (14087)
value ERROR_SXS_PROTECTION_CATALOG_FILE_MISSING (14078)
value ERROR_SXS_PROTECTION_CATALOG_NOT_VALID (14076)
value ERROR_SXS_PROTECTION_PUBLIC_KEY_TOO_SHORT (14075)
value ERROR_SXS_PROTECTION_RECOVERY_FAILED (14074)
value ERROR_SXS_RELEASE_ACTIVATION_CONTEXT (14088)
value ERROR_SXS_ROOT_MANIFEST_DEPENDENCY_NOT_INSTALLED (14015)
value ERROR_SXS_SECTION_NOT_FOUND (14000)
value ERROR_SXS_SETTING_NOT_REGISTERED (14106)
value ERROR_SXS_SYSTEM_DEFAULT_ACTIVATION_CONTEXT_EMPTY (14089)
value ERROR_SXS_THREAD_QUERIES_DISABLED (14010)
value ERROR_SXS_TRANSACTION_CLOSURE_INCOMPLETE (14107)
value ERROR_SXS_UNKNOWN_ENCODING (14013)
value ERROR_SXS_UNKNOWN_ENCODING_GROUP (14012)
value ERROR_SXS_UNTRANSLATABLE_HRESULT (14077)
value ERROR_SXS_VERSION_CONFLICT (14008)
value ERROR_SXS_WRONG_SECTION_TYPE (14009)
value ERROR_SXS_XML_E_BADCHARDATA (14036)
value ERROR_SXS_XML_E_BADCHARINSTRING (14034)
value ERROR_SXS_XML_E_BADNAMECHAR (14033)
value ERROR_SXS_XML_E_BADPEREFINSUBSET (14059)
value ERROR_SXS_XML_E_BADSTARTNAMECHAR (14032)
value ERROR_SXS_XML_E_BADXMLCASE (14069)
value ERROR_SXS_XML_E_BADXMLDECL (14056)
value ERROR_SXS_XML_E_COMMENTSYNTAX (14031)
value ERROR_SXS_XML_E_DUPLICATEATTRIBUTE (14053)
value ERROR_SXS_XML_E_EXPECTINGCLOSEQUOTE (14045)
value ERROR_SXS_XML_E_EXPECTINGTAGEND (14038)
value ERROR_SXS_XML_E_INCOMPLETE_ENCODING (14043)
value ERROR_SXS_XML_E_INTERNALERROR (14041)
value ERROR_SXS_XML_E_INVALIDATROOTLEVEL (14055)
value ERROR_SXS_XML_E_INVALIDENCODING (14067)
value ERROR_SXS_XML_E_INVALIDSWITCH (14068)
value ERROR_SXS_XML_E_INVALID_DECIMAL (14047)
value ERROR_SXS_XML_E_INVALID_HEXIDECIMAL (14048)
value ERROR_SXS_XML_E_INVALID_STANDALONE (14070)
value ERROR_SXS_XML_E_INVALID_UNICODE (14049)
value ERROR_SXS_XML_E_INVALID_VERSION (14072)
value ERROR_SXS_XML_E_MISSINGEQUALS (14073)
value ERROR_SXS_XML_E_MISSINGQUOTE (14030)
value ERROR_SXS_XML_E_MISSINGROOT (14057)
value ERROR_SXS_XML_E_MISSINGSEMICOLON (14039)
value ERROR_SXS_XML_E_MISSINGWHITESPACE (14037)
value ERROR_SXS_XML_E_MISSING_PAREN (14044)
value ERROR_SXS_XML_E_MULTIPLEROOTS (14054)
value ERROR_SXS_XML_E_MULTIPLE_COLONS (14046)
value ERROR_SXS_XML_E_RESERVEDNAMESPACE (14066)
value ERROR_SXS_XML_E_UNBALANCEDPAREN (14040)
value ERROR_SXS_XML_E_UNCLOSEDCDATA (14065)
value ERROR_SXS_XML_E_UNCLOSEDCOMMENT (14063)
value ERROR_SXS_XML_E_UNCLOSEDDECL (14064)
value ERROR_SXS_XML_E_UNCLOSEDENDTAG (14061)
value ERROR_SXS_XML_E_UNCLOSEDSTARTTAG (14060)
value ERROR_SXS_XML_E_UNCLOSEDSTRING (14062)
value ERROR_SXS_XML_E_UNCLOSEDTAG (14052)
value ERROR_SXS_XML_E_UNEXPECTEDENDTAG (14051)
value ERROR_SXS_XML_E_UNEXPECTEDEOF (14058)
value ERROR_SXS_XML_E_UNEXPECTED_STANDALONE (14071)
value ERROR_SXS_XML_E_UNEXPECTED_WHITESPACE (14042)
value ERROR_SXS_XML_E_WHITESPACEORQUESTIONMARK (14050)
value ERROR_SXS_XML_E_XMLDECLSYNTAX (14035)
value ERROR_SYMLINK_CLASS_DISABLED (1463)
value ERROR_SYMLINK_NOT_SUPPORTED (1464)
value ERROR_SYNCHRONIZATION_REQUIRED (569)
value ERROR_SYNC_FOREGROUND_REFRESH_REQUIRED (1274)
value ERROR_SYSTEM_DEVICE_NOT_FOUND (15299)
value ERROR_SYSTEM_HIVE_TOO_LARGE (653)
value ERROR_SYSTEM_IMAGE_BAD_SIGNATURE (637)
value ERROR_SYSTEM_INTEGRITY_INVALID_POLICY (4552)
value ERROR_SYSTEM_INTEGRITY_POLICY_NOT_SIGNED (4553)
value ERROR_SYSTEM_INTEGRITY_POLICY_VIOLATION (4551)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_DANGEROUS_EXT (4558)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_MALICIOUS (4556)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_OFFLINE (4559)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_PUA (4557)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_UNATTAINABLE (4581)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_UNFRIENDLY_FILE (4580)
value ERROR_SYSTEM_INTEGRITY_ROLLBACK_DETECTED (4550)
value ERROR_SYSTEM_INTEGRITY_SUPPLEMENTAL_POLICY_NOT_AUTHORIZED (4555)
value ERROR_SYSTEM_INTEGRITY_TOO_MANY_POLICIES (4554)
value ERROR_SYSTEM_NEEDS_REMEDIATION (15623)
value ERROR_SYSTEM_POWERSTATE_COMPLEX_TRANSITION (783)
value ERROR_SYSTEM_POWERSTATE_TRANSITION (782)
value ERROR_SYSTEM_PROCESS_TERMINATED (591)
value ERROR_SYSTEM_SHUTDOWN (641)
value ERROR_SYSTEM_TRACE (150)
value ERROR_TAG_NOT_FOUND (2012)
value ERROR_TAG_NOT_PRESENT (2013)
value ERROR_THREAD_ALREADY_IN_TASK (1552)
value ERROR_THREAD_MODE_ALREADY_BACKGROUND (400)
value ERROR_THREAD_MODE_NOT_BACKGROUND (401)
value ERROR_THREAD_NOT_IN_PROCESS (566)
value ERROR_THREAD_WAS_SUSPENDED (699)
value ERROR_TIERING_ALREADY_PROCESSING (_HRESULT_TYPEDEF_(0x80830006L))
value ERROR_TIERING_CANNOT_PIN_OBJECT (_HRESULT_TYPEDEF_(0x80830007L))
value ERROR_TIERING_FILE_IS_NOT_PINNED (_HRESULT_TYPEDEF_(0x80830008L))
value ERROR_TIERING_INVALID_FILE_ID (_HRESULT_TYPEDEF_(0x80830004L))
value ERROR_TIERING_NOT_SUPPORTED_ON_VOLUME (_HRESULT_TYPEDEF_(0x80830001L))
value ERROR_TIERING_STORAGE_TIER_NOT_FOUND (_HRESULT_TYPEDEF_(0x80830003L))
value ERROR_TIERING_VOLUME_DISMOUNT_IN_PROGRESS (_HRESULT_TYPEDEF_(0x80830002L))
value ERROR_TIERING_WRONG_CLUSTER_NODE (_HRESULT_TYPEDEF_(0x80830005L))
value ERROR_TIMEOUT (1460)
value ERROR_TIMER_NOT_CANCELED (541)
value ERROR_TIMER_RESOLUTION_NOT_SET (607)
value ERROR_TIMER_RESUME_IGNORED (722)
value ERROR_TIME_SENSITIVE_THREAD (422)
value ERROR_TIME_SKEW (1398)
value ERROR_TLW_WITH_WSCHILD (1406)
value ERROR_TM_IDENTITY_MISMATCH (6845)
value ERROR_TM_INITIALIZATION_FAILED (6706)
value ERROR_TM_VOLATILE (6828)
value ERROR_TOKEN_ALREADY_IN_USE (1375)
value ERROR_TOO_MANY_CMDS (56)
value ERROR_TOO_MANY_CONTEXT_IDS (1384)
value ERROR_TOO_MANY_DESCRIPTORS (331)
value ERROR_TOO_MANY_LINKS (1142)
value ERROR_TOO_MANY_LUIDS_REQUESTED (1333)
value ERROR_TOO_MANY_MODULES (214)
value ERROR_TOO_MANY_MUXWAITERS (152)
value ERROR_TOO_MANY_NAMES (68)
value ERROR_TOO_MANY_OPEN_FILES (4)
value ERROR_TOO_MANY_POSTS (298)
value ERROR_TOO_MANY_SECRETS (1381)
value ERROR_TOO_MANY_SEMAPHORES (100)
value ERROR_TOO_MANY_SEM_REQUESTS (103)
value ERROR_TOO_MANY_SESS (69)
value ERROR_TOO_MANY_SIDS (1389)
value ERROR_TOO_MANY_TCBS (155)
value ERROR_TOO_MANY_THREADS (565)
value ERROR_TRANSACTED_MAPPING_UNSUPPORTED_REMOTE (6834)
value ERROR_TRANSACTIONAL_CONFLICT (6800)
value ERROR_TRANSACTIONAL_OPEN_NOT_ALLOWED (6832)
value ERROR_TRANSACTIONMANAGER_IDENTITY_MISMATCH (6727)
value ERROR_TRANSACTIONMANAGER_NOT_FOUND (6718)
value ERROR_TRANSACTIONMANAGER_NOT_ONLINE (6719)
value ERROR_TRANSACTIONMANAGER_RECOVERY_NAME_COLLISION (6720)
value ERROR_TRANSACTIONS_NOT_FROZEN (6839)
value ERROR_TRANSACTIONS_UNSUPPORTED_REMOTE (6805)
value ERROR_TRANSACTION_ALREADY_ABORTED (6704)
value ERROR_TRANSACTION_ALREADY_COMMITTED (6705)
value ERROR_TRANSACTION_FREEZE_IN_PROGRESS (6840)
value ERROR_TRANSACTION_INTEGRITY_VIOLATED (6726)
value ERROR_TRANSACTION_INVALID_MARSHALL_BUFFER (6713)
value ERROR_TRANSACTION_MUST_WRITETHROUGH (6729)
value ERROR_TRANSACTION_NOT_ACTIVE (6701)
value ERROR_TRANSACTION_NOT_ENLISTED (6855)
value ERROR_TRANSACTION_NOT_FOUND (6715)
value ERROR_TRANSACTION_NOT_JOINED (6708)
value ERROR_TRANSACTION_NOT_REQUESTED (6703)
value ERROR_TRANSACTION_NOT_ROOT (6721)
value ERROR_TRANSACTION_NO_SUPERIOR (6730)
value ERROR_TRANSACTION_OBJECT_EXPIRED (6722)
value ERROR_TRANSACTION_PROPAGATION_FAILED (6711)
value ERROR_TRANSACTION_RECORD_TOO_LONG (6724)
value ERROR_TRANSACTION_REQUEST_NOT_VALID (6702)
value ERROR_TRANSACTION_REQUIRED_PROMOTION (6837)
value ERROR_TRANSACTION_RESPONSE_NOT_ENLISTED (6723)
value ERROR_TRANSACTION_SCOPE_CALLBACKS_NOT_SET (6836)
value ERROR_TRANSACTION_SUPERIOR_EXISTS (6709)
value ERROR_TRANSFORM_NOT_SUPPORTED (2004)
value ERROR_TRANSLATION_COMPLETE (757)
value ERROR_TRANSPORT_FULL (4328)
value ERROR_TRAY_MALFUNCTION (0x00000010)
value ERROR_TRUSTED_DOMAIN_FAILURE (1788)
value ERROR_TRUSTED_RELATIONSHIP_FAILURE (1789)
value ERROR_TRUST_FAILURE (1790)
value ERROR_TS_INCOMPATIBLE_SESSIONS (7069)
value ERROR_TS_VIDEO_SUBSYSTEM_ERROR (7070)
value ERROR_TXF_ATTRIBUTE_CORRUPT (6830)
value ERROR_TXF_DIR_NOT_EMPTY (6826)
value ERROR_TXF_METADATA_ALREADY_PRESENT (6835)
value ERROR_UNABLE_TO_CLEAN (4311)
value ERROR_UNABLE_TO_EJECT_MOUNTED_MEDIA (4330)
value ERROR_UNABLE_TO_INVENTORY_DRIVE (4325)
value ERROR_UNABLE_TO_INVENTORY_SLOT (4326)
value ERROR_UNABLE_TO_INVENTORY_TRANSPORT (4327)
value ERROR_UNABLE_TO_LOAD_MEDIUM (4324)
value ERROR_UNABLE_TO_LOCK_MEDIA (1108)
value ERROR_UNABLE_TO_MOVE_REPLACEMENT (1176)
value ERROR_UNABLE_TO_REMOVE_REPLACED (1175)
value ERROR_UNABLE_TO_UNLOAD_MEDIA (1109)
value ERROR_UNDEFINED_CHARACTER (583)
value ERROR_UNDEFINED_SCOPE (319)
value ERROR_UNEXPECTED_MM_CREATE_ERR (556)
value ERROR_UNEXPECTED_MM_EXTEND_ERR (558)
value ERROR_UNEXPECTED_MM_MAP_ERROR (557)
value ERROR_UNEXPECTED_NTCACHEMANAGER_ERROR (443)
value ERROR_UNEXPECTED_OMID (4334)
value ERROR_UNEXP_NET_ERR (59)
value ERROR_UNHANDLED_ERROR (0xFFFFFFFF)
value ERROR_UNHANDLED_EXCEPTION (574)
value ERROR_UNIDENTIFIED_ERROR (1287)
value ERROR_UNKNOWN_COMPONENT (1607)
value ERROR_UNKNOWN_FEATURE (1606)
value ERROR_UNKNOWN_PATCH (1647)
value ERROR_UNKNOWN_PORT (1796)
value ERROR_UNKNOWN_PRINTER_DRIVER (1797)
value ERROR_UNKNOWN_PRINTPROCESSOR (1798)
value ERROR_UNKNOWN_PRINT_MONITOR (3000)
value ERROR_UNKNOWN_PRODUCT (1605)
value ERROR_UNKNOWN_PROPERTY (1608)
value ERROR_UNKNOWN_REVISION (1305)
value ERROR_UNMAPPED_SUBSTITUTION_STRING (14096)
value ERROR_UNRECOGNIZED_MEDIA (1785)
value ERROR_UNRECOGNIZED_VOLUME (1005)
value ERROR_UNSATISFIED_DEPENDENCIES (441)
value ERROR_UNSIGNED_PACKAGE_INVALID_CONTENT (15659)
value ERROR_UNSIGNED_PACKAGE_INVALID_PUBLISHER_NAMESPACE (15660)
value ERROR_UNSUPPORTED_COMPRESSION (618)
value ERROR_UNSUPPORTED_TYPE (1630)
value ERROR_UNTRUSTED_MOUNT_POINT (448)
value ERROR_UNWIND (542)
value ERROR_UNWIND_CONSOLIDATE (684)
value ERROR_USER_APC (737)
value ERROR_USER_DELETE_TRUST_QUOTA_EXCEEDED (1934)
value ERROR_USER_EXISTS (1316)
value ERROR_USER_MAPPED_FILE (1224)
value ERROR_USER_PROFILE_LOAD (500)
value ERROR_VALIDATE_CONTINUE (625)
value ERROR_VC_DISCONNECTED (240)
value ERROR_VDM_DISALLOWED (1286)
value ERROR_VDM_HARD_ERROR (593)
value ERROR_VERIFIER_STOP (537)
value ERROR_VERSION_PARSE_ERROR (777)
value ERROR_VHDSET_BACKING_STORAGE_NOT_FOUND (_HRESULT_TYPEDEF_(0xC05CFF0CL))
value ERROR_VHD_ALREADY_AT_OR_BELOW_MINIMUM_VIRTUAL_SIZE (_NDIS_ERROR_TYPEDEF_(0xC03A0027L))
value ERROR_VHD_BITMAP_MISMATCH (_NDIS_ERROR_TYPEDEF_(0xC03A000CL))
value ERROR_VHD_BLOCK_ALLOCATION_FAILURE (_NDIS_ERROR_TYPEDEF_(0xC03A0009L))
value ERROR_VHD_BLOCK_ALLOCATION_TABLE_CORRUPT (_NDIS_ERROR_TYPEDEF_(0xC03A000AL))
value ERROR_VHD_CHANGE_TRACKING_DISABLED (_NDIS_ERROR_TYPEDEF_(0xC03A002AL))
value ERROR_VHD_CHILD_PARENT_ID_MISMATCH (_NDIS_ERROR_TYPEDEF_(0xC03A000EL))
value ERROR_VHD_CHILD_PARENT_SIZE_MISMATCH (_NDIS_ERROR_TYPEDEF_(0xC03A0017L))
value ERROR_VHD_CHILD_PARENT_TIMESTAMP_MISMATCH (_NDIS_ERROR_TYPEDEF_(0xC03A000FL))
value ERROR_VHD_COULD_NOT_COMPUTE_MINIMUM_VIRTUAL_SIZE (_NDIS_ERROR_TYPEDEF_(0xC03A0026L))
value ERROR_VHD_DIFFERENCING_CHAIN_CYCLE_DETECTED (_NDIS_ERROR_TYPEDEF_(0xC03A0018L))
value ERROR_VHD_DIFFERENCING_CHAIN_ERROR_IN_PARENT (_NDIS_ERROR_TYPEDEF_(0xC03A0019L))
value ERROR_VHD_DRIVE_FOOTER_CHECKSUM_MISMATCH (_NDIS_ERROR_TYPEDEF_(0xC03A0002L))
value ERROR_VHD_DRIVE_FOOTER_CORRUPT (_NDIS_ERROR_TYPEDEF_(0xC03A0003L))
value ERROR_VHD_DRIVE_FOOTER_MISSING (_NDIS_ERROR_TYPEDEF_(0xC03A0001L))
value ERROR_VHD_FORMAT_UNKNOWN (_NDIS_ERROR_TYPEDEF_(0xC03A0004L))
value ERROR_VHD_FORMAT_UNSUPPORTED_VERSION (_NDIS_ERROR_TYPEDEF_(0xC03A0005L))
value ERROR_VHD_INVALID_BLOCK_SIZE (_NDIS_ERROR_TYPEDEF_(0xC03A000BL))
value ERROR_VHD_INVALID_CHANGE_TRACKING_ID (_NDIS_ERROR_TYPEDEF_(0xC03A0029L))
value ERROR_VHD_INVALID_FILE_SIZE (_NDIS_ERROR_TYPEDEF_(0xC03A0013L))
value ERROR_VHD_INVALID_SIZE (_NDIS_ERROR_TYPEDEF_(0xC03A0012L))
value ERROR_VHD_INVALID_STATE (_NDIS_ERROR_TYPEDEF_(0xC03A001CL))
value ERROR_VHD_INVALID_TYPE (_NDIS_ERROR_TYPEDEF_(0xC03A001BL))
value ERROR_VHD_METADATA_FULL (_NDIS_ERROR_TYPEDEF_(0xC03A0028L))
value ERROR_VHD_METADATA_READ_FAILURE (_NDIS_ERROR_TYPEDEF_(0xC03A0010L))
value ERROR_VHD_METADATA_WRITE_FAILURE (_NDIS_ERROR_TYPEDEF_(0xC03A0011L))
value ERROR_VHD_MISSING_CHANGE_TRACKING_INFORMATION (_NDIS_ERROR_TYPEDEF_(0xC03A0030L))
value ERROR_VHD_PARENT_VHD_ACCESS_DENIED (_NDIS_ERROR_TYPEDEF_(0xC03A0016L))
value ERROR_VHD_PARENT_VHD_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0xC03A000DL))
value ERROR_VHD_RESIZE_WOULD_TRUNCATE_DATA (_NDIS_ERROR_TYPEDEF_(0xC03A0025L))
value ERROR_VHD_SHARED (_HRESULT_TYPEDEF_(0xC05CFF0AL))
value ERROR_VHD_SPARSE_HEADER_CHECKSUM_MISMATCH (_NDIS_ERROR_TYPEDEF_(0xC03A0006L))
value ERROR_VHD_SPARSE_HEADER_CORRUPT (_NDIS_ERROR_TYPEDEF_(0xC03A0008L))
value ERROR_VHD_SPARSE_HEADER_UNSUPPORTED_VERSION (_NDIS_ERROR_TYPEDEF_(0xC03A0007L))
value ERROR_VID_CHILD_GPA_PAGE_SET_CORRUPTED (_NDIS_ERROR_TYPEDEF_(0xC037000EL))
value ERROR_VID_DUPLICATE_HANDLER (_NDIS_ERROR_TYPEDEF_(0xC0370001L))
value ERROR_VID_EXCEEDED_KM_CONTEXT_COUNT_LIMIT (_NDIS_ERROR_TYPEDEF_(0xC037001EL))
value ERROR_VID_EXCEEDED_MBP_ENTRY_MAP_LIMIT (_NDIS_ERROR_TYPEDEF_(0xC037000CL))
value ERROR_VID_HANDLER_NOT_PRESENT (_NDIS_ERROR_TYPEDEF_(0xC0370004L))
value ERROR_VID_INSUFFICIENT_RESOURCES_HV_DEPOSIT (_NDIS_ERROR_TYPEDEF_(0xC037002DL))
value ERROR_VID_INSUFFICIENT_RESOURCES_PHYSICAL_BUFFER (_NDIS_ERROR_TYPEDEF_(0xC037002CL))
value ERROR_VID_INSUFFICIENT_RESOURCES_RESERVE (_NDIS_ERROR_TYPEDEF_(0xC037002BL))
value ERROR_VID_INSUFFICIENT_RESOURCES_WITHDRAW (_NDIS_ERROR_TYPEDEF_(0xC037002FL))
value ERROR_VID_INVALID_CHILD_GPA_PAGE_SET (_NDIS_ERROR_TYPEDEF_(0xC0370022L))
value ERROR_VID_INVALID_GPA_RANGE_HANDLE (_NDIS_ERROR_TYPEDEF_(0xC0370015L))
value ERROR_VID_INVALID_MEMORY_BLOCK_HANDLE (_NDIS_ERROR_TYPEDEF_(0xC0370012L))
value ERROR_VID_INVALID_MESSAGE_QUEUE_HANDLE (_NDIS_ERROR_TYPEDEF_(0xC0370014L))
value ERROR_VID_INVALID_NUMA_NODE_INDEX (_NDIS_ERROR_TYPEDEF_(0xC0370010L))
value ERROR_VID_INVALID_NUMA_SETTINGS (_NDIS_ERROR_TYPEDEF_(0xC037000FL))
value ERROR_VID_INVALID_OBJECT_NAME (_NDIS_ERROR_TYPEDEF_(0xC0370005L))
value ERROR_VID_INVALID_PPM_HANDLE (_NDIS_ERROR_TYPEDEF_(0xC0370018L))
value ERROR_VID_INVALID_PROCESSOR_STATE (_NDIS_ERROR_TYPEDEF_(0xC037001DL))
value ERROR_VID_KM_INTERFACE_ALREADY_INITIALIZED (_NDIS_ERROR_TYPEDEF_(0xC037001FL))
value ERROR_VID_MBPS_ARE_LOCKED (_NDIS_ERROR_TYPEDEF_(0xC0370019L))
value ERROR_VID_MBP_ALREADY_LOCKED_USING_RESERVED_PAGE (_NDIS_ERROR_TYPEDEF_(0xC0370025L))
value ERROR_VID_MBP_COUNT_EXCEEDED_LIMIT (_NDIS_ERROR_TYPEDEF_(0xC0370026L))
value ERROR_VID_MB_PROPERTY_ALREADY_SET_RESET (_NDIS_ERROR_TYPEDEF_(0xC0370020L))
value ERROR_VID_MB_STILL_REFERENCED (_NDIS_ERROR_TYPEDEF_(0xC037000DL))
value ERROR_VID_MEMORY_BLOCK_LOCK_COUNT_EXCEEDED (_NDIS_ERROR_TYPEDEF_(0xC0370017L))
value ERROR_VID_MEMORY_TYPE_NOT_SUPPORTED (_NDIS_ERROR_TYPEDEF_(0xC037002EL))
value ERROR_VID_MESSAGE_QUEUE_ALREADY_EXISTS (_NDIS_ERROR_TYPEDEF_(0xC037000BL))
value ERROR_VID_MESSAGE_QUEUE_CLOSED (_NDIS_ERROR_TYPEDEF_(0xC037001AL))
value ERROR_VID_MESSAGE_QUEUE_NAME_TOO_LONG (_NDIS_ERROR_TYPEDEF_(0xC0370007L))
value ERROR_VID_MMIO_RANGE_DESTROYED (_NDIS_ERROR_TYPEDEF_(0xC0370021L))
value ERROR_VID_NOTIFICATION_QUEUE_ALREADY_ASSOCIATED (_NDIS_ERROR_TYPEDEF_(0xC0370011L))
value ERROR_VID_NO_MEMORY_BLOCK_NOTIFICATION_QUEUE (_NDIS_ERROR_TYPEDEF_(0xC0370016L))
value ERROR_VID_PAGE_RANGE_OVERFLOW (_NDIS_ERROR_TYPEDEF_(0xC0370013L))
value ERROR_VID_PARTITION_ALREADY_EXISTS (_NDIS_ERROR_TYPEDEF_(0xC0370008L))
value ERROR_VID_PARTITION_DOES_NOT_EXIST (_NDIS_ERROR_TYPEDEF_(0xC0370009L))
value ERROR_VID_PARTITION_NAME_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0xC037000AL))
value ERROR_VID_PARTITION_NAME_TOO_LONG (_NDIS_ERROR_TYPEDEF_(0xC0370006L))
value ERROR_VID_PROCESS_ALREADY_SET (_NDIS_ERROR_TYPEDEF_(0xC0370030L))
value ERROR_VID_QUEUE_FULL (_NDIS_ERROR_TYPEDEF_(0xC0370003L))
value ERROR_VID_REMOTE_NODE_PARENT_GPA_PAGES_USED (_NDIS_ERROR_TYPEDEF_(0x80370001L))
value ERROR_VID_RESERVE_PAGE_SET_IS_BEING_USED (_NDIS_ERROR_TYPEDEF_(0xC0370023L))
value ERROR_VID_RESERVE_PAGE_SET_TOO_SMALL (_NDIS_ERROR_TYPEDEF_(0xC0370024L))
value ERROR_VID_SAVED_STATE_CORRUPT (_NDIS_ERROR_TYPEDEF_(0xC0370027L))
value ERROR_VID_SAVED_STATE_INCOMPATIBLE (_NDIS_ERROR_TYPEDEF_(0xC0370029L))
value ERROR_VID_SAVED_STATE_UNRECOGNIZED_ITEM (_NDIS_ERROR_TYPEDEF_(0xC0370028L))
value ERROR_VID_STOP_PENDING (_NDIS_ERROR_TYPEDEF_(0xC037001CL))
value ERROR_VID_TOO_MANY_HANDLERS (_NDIS_ERROR_TYPEDEF_(0xC0370002L))
value ERROR_VID_VIRTUAL_PROCESSOR_LIMIT_EXCEEDED (_NDIS_ERROR_TYPEDEF_(0xC037001BL))
value ERROR_VID_VTL_ACCESS_DENIED (_NDIS_ERROR_TYPEDEF_(0xC037002AL))
value ERROR_VIRTDISK_DISK_ALREADY_OWNED (_NDIS_ERROR_TYPEDEF_(0xC03A001EL))
value ERROR_VIRTDISK_DISK_ONLINE_AND_WRITABLE (_NDIS_ERROR_TYPEDEF_(0xC03A001FL))
value ERROR_VIRTDISK_NOT_VIRTUAL_DISK (_NDIS_ERROR_TYPEDEF_(0xC03A0015L))
value ERROR_VIRTDISK_PROVIDER_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0xC03A0014L))
value ERROR_VIRTDISK_UNSUPPORTED_DISK_SECTOR_SIZE (_NDIS_ERROR_TYPEDEF_(0xC03A001DL))
value ERROR_VIRTUAL_DISK_LIMITATION (_NDIS_ERROR_TYPEDEF_(0xC03A001AL))
value ERROR_VIRUS_DELETED (226)
value ERROR_VIRUS_INFECTED (225)
value ERROR_VMCOMPUTE_CONNECTION_CLOSED (_NDIS_ERROR_TYPEDEF_(0xC037010AL))
value ERROR_VMCOMPUTE_CONNECT_FAILED (_NDIS_ERROR_TYPEDEF_(0xC0370108L))
value ERROR_VMCOMPUTE_HYPERV_NOT_INSTALLED (_NDIS_ERROR_TYPEDEF_(0xC0370102L))
value ERROR_VMCOMPUTE_IMAGE_MISMATCH (_NDIS_ERROR_TYPEDEF_(0xC0370101L))
value ERROR_VMCOMPUTE_INVALID_JSON (_NDIS_ERROR_TYPEDEF_(0xC037010DL))
value ERROR_VMCOMPUTE_INVALID_LAYER (_NDIS_ERROR_TYPEDEF_(0xC0370112L))
value ERROR_VMCOMPUTE_INVALID_STATE (_NDIS_ERROR_TYPEDEF_(0xC0370105L))
value ERROR_VMCOMPUTE_OPERATION_PENDING (_NDIS_ERROR_TYPEDEF_(0xC0370103L))
value ERROR_VMCOMPUTE_PROTOCOL_ERROR (_NDIS_ERROR_TYPEDEF_(0xC0370111L))
value ERROR_VMCOMPUTE_SYSTEM_ALREADY_EXISTS (_NDIS_ERROR_TYPEDEF_(0xC037010FL))
value ERROR_VMCOMPUTE_SYSTEM_ALREADY_STOPPED (_NDIS_ERROR_TYPEDEF_(0xC0370110L))
value ERROR_VMCOMPUTE_SYSTEM_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0xC037010EL))
value ERROR_VMCOMPUTE_TERMINATED (_NDIS_ERROR_TYPEDEF_(0xC0370107L))
value ERROR_VMCOMPUTE_TERMINATED_DURING_START (_NDIS_ERROR_TYPEDEF_(0xC0370100L))
value ERROR_VMCOMPUTE_TIMEOUT (_NDIS_ERROR_TYPEDEF_(0xC0370109L))
value ERROR_VMCOMPUTE_TOO_MANY_NOTIFICATIONS (_NDIS_ERROR_TYPEDEF_(0xC0370104L))
value ERROR_VMCOMPUTE_UNEXPECTED_EXIT (_NDIS_ERROR_TYPEDEF_(0xC0370106L))
value ERROR_VMCOMPUTE_UNKNOWN_MESSAGE (_NDIS_ERROR_TYPEDEF_(0xC037010BL))
value ERROR_VMCOMPUTE_UNSUPPORTED_PROTOCOL_VERSION (_NDIS_ERROR_TYPEDEF_(0xC037010CL))
value ERROR_VMCOMPUTE_WINDOWS_INSIDER_REQUIRED (_NDIS_ERROR_TYPEDEF_(0xC0370113L))
value ERROR_VNET_VIRTUAL_SWITCH_NAME_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0xC0370200L))
value ERROR_VOLMGR_ALL_DISKS_FAILED (_NDIS_ERROR_TYPEDEF_(0xC0380029L))
value ERROR_VOLMGR_BAD_BOOT_DISK (_NDIS_ERROR_TYPEDEF_(0xC038004FL))
value ERROR_VOLMGR_DATABASE_FULL (_NDIS_ERROR_TYPEDEF_(0xC0380001L))
value ERROR_VOLMGR_DIFFERENT_SECTOR_SIZE (_NDIS_ERROR_TYPEDEF_(0xC038004EL))
value ERROR_VOLMGR_DISK_CONFIGURATION_CORRUPTED (_NDIS_ERROR_TYPEDEF_(0xC0380002L))
value ERROR_VOLMGR_DISK_CONFIGURATION_NOT_IN_SYNC (_NDIS_ERROR_TYPEDEF_(0xC0380003L))
value ERROR_VOLMGR_DISK_CONTAINS_NON_SIMPLE_VOLUME (_NDIS_ERROR_TYPEDEF_(0xC0380005L))
value ERROR_VOLMGR_DISK_DUPLICATE (_NDIS_ERROR_TYPEDEF_(0xC0380006L))
value ERROR_VOLMGR_DISK_DYNAMIC (_NDIS_ERROR_TYPEDEF_(0xC0380007L))
value ERROR_VOLMGR_DISK_ID_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380008L))
value ERROR_VOLMGR_DISK_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380009L))
value ERROR_VOLMGR_DISK_LAST_VOTER (_NDIS_ERROR_TYPEDEF_(0xC038000AL))
value ERROR_VOLMGR_DISK_LAYOUT_INVALID (_NDIS_ERROR_TYPEDEF_(0xC038000BL))
value ERROR_VOLMGR_DISK_LAYOUT_NON_BASIC_BETWEEN_BASIC_PARTITIONS (_NDIS_ERROR_TYPEDEF_(0xC038000CL))
value ERROR_VOLMGR_DISK_LAYOUT_NOT_CYLINDER_ALIGNED (_NDIS_ERROR_TYPEDEF_(0xC038000DL))
value ERROR_VOLMGR_DISK_LAYOUT_PARTITIONS_TOO_SMALL (_NDIS_ERROR_TYPEDEF_(0xC038000EL))
value ERROR_VOLMGR_DISK_LAYOUT_PRIMARY_BETWEEN_LOGICAL_PARTITIONS (_NDIS_ERROR_TYPEDEF_(0xC038000FL))
value ERROR_VOLMGR_DISK_LAYOUT_TOO_MANY_PARTITIONS (_NDIS_ERROR_TYPEDEF_(0xC0380010L))
value ERROR_VOLMGR_DISK_MISSING (_NDIS_ERROR_TYPEDEF_(0xC0380011L))
value ERROR_VOLMGR_DISK_NOT_EMPTY (_NDIS_ERROR_TYPEDEF_(0xC0380012L))
value ERROR_VOLMGR_DISK_NOT_ENOUGH_SPACE (_NDIS_ERROR_TYPEDEF_(0xC0380013L))
value ERROR_VOLMGR_DISK_REVECTORING_FAILED (_NDIS_ERROR_TYPEDEF_(0xC0380014L))
value ERROR_VOLMGR_DISK_SECTOR_SIZE_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380015L))
value ERROR_VOLMGR_DISK_SET_NOT_CONTAINED (_NDIS_ERROR_TYPEDEF_(0xC0380016L))
value ERROR_VOLMGR_DISK_USED_BY_MULTIPLE_MEMBERS (_NDIS_ERROR_TYPEDEF_(0xC0380017L))
value ERROR_VOLMGR_DISK_USED_BY_MULTIPLE_PLEXES (_NDIS_ERROR_TYPEDEF_(0xC0380018L))
value ERROR_VOLMGR_DYNAMIC_DISK_NOT_SUPPORTED (_NDIS_ERROR_TYPEDEF_(0xC0380019L))
value ERROR_VOLMGR_EXTENT_ALREADY_USED (_NDIS_ERROR_TYPEDEF_(0xC038001AL))
value ERROR_VOLMGR_EXTENT_NOT_CONTIGUOUS (_NDIS_ERROR_TYPEDEF_(0xC038001BL))
value ERROR_VOLMGR_EXTENT_NOT_IN_PUBLIC_REGION (_NDIS_ERROR_TYPEDEF_(0xC038001CL))
value ERROR_VOLMGR_EXTENT_NOT_SECTOR_ALIGNED (_NDIS_ERROR_TYPEDEF_(0xC038001DL))
value ERROR_VOLMGR_EXTENT_OVERLAPS_EBR_PARTITION (_NDIS_ERROR_TYPEDEF_(0xC038001EL))
value ERROR_VOLMGR_EXTENT_VOLUME_LENGTHS_DO_NOT_MATCH (_NDIS_ERROR_TYPEDEF_(0xC038001FL))
value ERROR_VOLMGR_FAULT_TOLERANT_NOT_SUPPORTED (_NDIS_ERROR_TYPEDEF_(0xC0380020L))
value ERROR_VOLMGR_INCOMPLETE_DISK_MIGRATION (_NDIS_ERROR_TYPEDEF_(0x80380002L))
value ERROR_VOLMGR_INCOMPLETE_REGENERATION (_NDIS_ERROR_TYPEDEF_(0x80380001L))
value ERROR_VOLMGR_INTERLEAVE_LENGTH_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380021L))
value ERROR_VOLMGR_MAXIMUM_REGISTERED_USERS (_NDIS_ERROR_TYPEDEF_(0xC0380022L))
value ERROR_VOLMGR_MEMBER_INDEX_DUPLICATE (_NDIS_ERROR_TYPEDEF_(0xC0380024L))
value ERROR_VOLMGR_MEMBER_INDEX_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380025L))
value ERROR_VOLMGR_MEMBER_IN_SYNC (_NDIS_ERROR_TYPEDEF_(0xC0380023L))
value ERROR_VOLMGR_MEMBER_MISSING (_NDIS_ERROR_TYPEDEF_(0xC0380026L))
value ERROR_VOLMGR_MEMBER_NOT_DETACHED (_NDIS_ERROR_TYPEDEF_(0xC0380027L))
value ERROR_VOLMGR_MEMBER_REGENERATING (_NDIS_ERROR_TYPEDEF_(0xC0380028L))
value ERROR_VOLMGR_MIRROR_NOT_SUPPORTED (_NDIS_ERROR_TYPEDEF_(0xC038005BL))
value ERROR_VOLMGR_NOTIFICATION_RESET (_NDIS_ERROR_TYPEDEF_(0xC038002CL))
value ERROR_VOLMGR_NOT_PRIMARY_PACK (_NDIS_ERROR_TYPEDEF_(0xC0380052L))
value ERROR_VOLMGR_NO_REGISTERED_USERS (_NDIS_ERROR_TYPEDEF_(0xC038002AL))
value ERROR_VOLMGR_NO_SUCH_USER (_NDIS_ERROR_TYPEDEF_(0xC038002BL))
value ERROR_VOLMGR_NO_VALID_LOG_COPIES (_NDIS_ERROR_TYPEDEF_(0xC0380058L))
value ERROR_VOLMGR_NUMBER_OF_DISKS_INVALID (_NDIS_ERROR_TYPEDEF_(0xC038005AL))
value ERROR_VOLMGR_NUMBER_OF_DISKS_IN_MEMBER_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380055L))
value ERROR_VOLMGR_NUMBER_OF_DISKS_IN_PLEX_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380054L))
value ERROR_VOLMGR_NUMBER_OF_EXTENTS_INVALID (_NDIS_ERROR_TYPEDEF_(0xC038004DL))
value ERROR_VOLMGR_NUMBER_OF_MEMBERS_INVALID (_NDIS_ERROR_TYPEDEF_(0xC038002DL))
value ERROR_VOLMGR_NUMBER_OF_PLEXES_INVALID (_NDIS_ERROR_TYPEDEF_(0xC038002EL))
value ERROR_VOLMGR_PACK_CONFIG_OFFLINE (_NDIS_ERROR_TYPEDEF_(0xC0380050L))
value ERROR_VOLMGR_PACK_CONFIG_ONLINE (_NDIS_ERROR_TYPEDEF_(0xC0380051L))
value ERROR_VOLMGR_PACK_CONFIG_UPDATE_FAILED (_NDIS_ERROR_TYPEDEF_(0xC0380004L))
value ERROR_VOLMGR_PACK_DUPLICATE (_NDIS_ERROR_TYPEDEF_(0xC038002FL))
value ERROR_VOLMGR_PACK_HAS_QUORUM (_NDIS_ERROR_TYPEDEF_(0xC0380034L))
value ERROR_VOLMGR_PACK_ID_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380030L))
value ERROR_VOLMGR_PACK_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380031L))
value ERROR_VOLMGR_PACK_LOG_UPDATE_FAILED (_NDIS_ERROR_TYPEDEF_(0xC0380053L))
value ERROR_VOLMGR_PACK_NAME_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380032L))
value ERROR_VOLMGR_PACK_OFFLINE (_NDIS_ERROR_TYPEDEF_(0xC0380033L))
value ERROR_VOLMGR_PACK_WITHOUT_QUORUM (_NDIS_ERROR_TYPEDEF_(0xC0380035L))
value ERROR_VOLMGR_PARTITION_STYLE_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380036L))
value ERROR_VOLMGR_PARTITION_UPDATE_FAILED (_NDIS_ERROR_TYPEDEF_(0xC0380037L))
value ERROR_VOLMGR_PLEX_INDEX_DUPLICATE (_NDIS_ERROR_TYPEDEF_(0xC0380039L))
value ERROR_VOLMGR_PLEX_INDEX_INVALID (_NDIS_ERROR_TYPEDEF_(0xC038003AL))
value ERROR_VOLMGR_PLEX_IN_SYNC (_NDIS_ERROR_TYPEDEF_(0xC0380038L))
value ERROR_VOLMGR_PLEX_LAST_ACTIVE (_NDIS_ERROR_TYPEDEF_(0xC038003BL))
value ERROR_VOLMGR_PLEX_MISSING (_NDIS_ERROR_TYPEDEF_(0xC038003CL))
value ERROR_VOLMGR_PLEX_NOT_SIMPLE (_NDIS_ERROR_TYPEDEF_(0xC0380040L))
value ERROR_VOLMGR_PLEX_NOT_SIMPLE_SPANNED (_NDIS_ERROR_TYPEDEF_(0xC0380057L))
value ERROR_VOLMGR_PLEX_REGENERATING (_NDIS_ERROR_TYPEDEF_(0xC038003DL))
value ERROR_VOLMGR_PLEX_TYPE_INVALID (_NDIS_ERROR_TYPEDEF_(0xC038003EL))
value ERROR_VOLMGR_PRIMARY_PACK_PRESENT (_NDIS_ERROR_TYPEDEF_(0xC0380059L))
value ERROR_VOLMGR_STRUCTURE_SIZE_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380041L))
value ERROR_VOLMGR_TOO_MANY_NOTIFICATION_REQUESTS (_NDIS_ERROR_TYPEDEF_(0xC0380042L))
value ERROR_VOLMGR_TRANSACTION_IN_PROGRESS (_NDIS_ERROR_TYPEDEF_(0xC0380043L))
value ERROR_VOLMGR_UNEXPECTED_DISK_LAYOUT_CHANGE (_NDIS_ERROR_TYPEDEF_(0xC0380044L))
value ERROR_VOLMGR_VOLUME_CONTAINS_MISSING_DISK (_NDIS_ERROR_TYPEDEF_(0xC0380045L))
value ERROR_VOLMGR_VOLUME_ID_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380046L))
value ERROR_VOLMGR_VOLUME_LENGTH_INVALID (_NDIS_ERROR_TYPEDEF_(0xC0380047L))
value ERROR_VOLMGR_VOLUME_LENGTH_NOT_SECTOR_SIZE_MULTIPLE (_NDIS_ERROR_TYPEDEF_(0xC0380048L))
value ERROR_VOLMGR_VOLUME_MIRRORED (_NDIS_ERROR_TYPEDEF_(0xC0380056L))
value ERROR_VOLMGR_VOLUME_NOT_MIRRORED (_NDIS_ERROR_TYPEDEF_(0xC0380049L))
value ERROR_VOLMGR_VOLUME_NOT_RETAINED (_NDIS_ERROR_TYPEDEF_(0xC038004AL))
value ERROR_VOLMGR_VOLUME_OFFLINE (_NDIS_ERROR_TYPEDEF_(0xC038004BL))
value ERROR_VOLMGR_VOLUME_RETAINED (_NDIS_ERROR_TYPEDEF_(0xC038004CL))
value ERROR_VOLSNAP_ACTIVATION_TIMEOUT (_HRESULT_TYPEDEF_(0x80820002L))
value ERROR_VOLSNAP_BOOTFILE_NOT_VALID (_HRESULT_TYPEDEF_(0x80820001L))
value ERROR_VOLSNAP_HIBERNATE_READY (761)
value ERROR_VOLSNAP_NO_BYPASSIO_WITH_SNAPSHOT (_HRESULT_TYPEDEF_(0x80820003L))
value ERROR_VOLSNAP_PREPARE_HIBERNATE (655)
value ERROR_VOLUME_CONTAINS_SYS_FILES (4337)
value ERROR_VOLUME_DIRTY (6851)
value ERROR_VOLUME_MOUNTED (743)
value ERROR_VOLUME_NOT_CLUSTER_ALIGNED (407)
value ERROR_VOLUME_NOT_SIS_ENABLED (4500)
value ERROR_VOLUME_NOT_SUPPORTED (492)
value ERROR_VOLUME_NOT_SUPPORT_EFS (6014)
value ERROR_VOLUME_WRITE_ACCESS_DENIED (508)
value ERROR_VRF_VOLATILE_CFG_AND_IO_ENABLED (3080)
value ERROR_VRF_VOLATILE_NMI_REGISTERED (3086)
value ERROR_VRF_VOLATILE_NOT_RUNNABLE_SYSTEM (3083)
value ERROR_VRF_VOLATILE_NOT_STOPPABLE (3081)
value ERROR_VRF_VOLATILE_NOT_SUPPORTED_RULECLASS (3084)
value ERROR_VRF_VOLATILE_PROTECTED_DRIVER (3085)
value ERROR_VRF_VOLATILE_SAFE_MODE (3082)
value ERROR_VRF_VOLATILE_SETTINGS_CONFLICT (3087)
value ERROR_VSMB_SAVED_STATE_CORRUPT (_NDIS_ERROR_TYPEDEF_(0xC0370401L))
value ERROR_VSMB_SAVED_STATE_FILE_NOT_FOUND (_NDIS_ERROR_TYPEDEF_(0xC0370400L))
value ERROR_VSM_DMA_PROTECTION_NOT_IN_USE (4561)
value ERROR_VSM_NOT_INITIALIZED (4560)
value ERROR_WAIT_FOR_OPLOCK (765)
value ERROR_WAIT_NO_CHILDREN (128)
value ERROR_WAKE_SYSTEM (730)
value ERROR_WAKE_SYSTEM_DEBUGGER (675)
value ERROR_WAS_LOCKED (717)
value ERROR_WAS_UNLOCKED (715)
value ERROR_WEAK_WHFBKEY_BLOCKED (8651)
value ERROR_WINDOW_NOT_COMBOBOX (1423)
value ERROR_WINDOW_NOT_DIALOG (1420)
value ERROR_WINDOW_OF_OTHER_THREAD (1408)
value ERROR_WINS_INTERNAL (4000)
value ERROR_WIP_ENCRYPTION_FAILED (6023)
value ERROR_WMI_ALREADY_DISABLED (4212)
value ERROR_WMI_ALREADY_ENABLED (4206)
value ERROR_WMI_DP_FAILED (4209)
value ERROR_WMI_DP_NOT_FOUND (4204)
value ERROR_WMI_GUID_DISCONNECTED (4207)
value ERROR_WMI_GUID_NOT_FOUND (4200)
value ERROR_WMI_INSTANCE_NOT_FOUND (4201)
value ERROR_WMI_INVALID_MOF (4210)
value ERROR_WMI_INVALID_REGINFO (4211)
value ERROR_WMI_ITEMID_NOT_FOUND (4202)
value ERROR_WMI_READ_ONLY (4213)
value ERROR_WMI_SERVER_UNAVAILABLE (4208)
value ERROR_WMI_SET_FAILURE (4214)
value ERROR_WMI_TRY_AGAIN (4203)
value ERROR_WMI_UNRESOLVED_INSTANCE_REF (4205)
value ERROR_WOF_FILE_RESOURCE_TABLE_CORRUPT (4448)
value ERROR_WOF_WIM_HEADER_CORRUPT (4446)
value ERROR_WOF_WIM_RESOURCE_TABLE_CORRUPT (4447)
value ERROR_WORKING_SET_QUOTA (1453)
value ERROR_WOW_ASSERTION (670)
value ERROR_WRITE_FAULT (29)
value ERROR_WRITE_PROTECT (19)
value ERROR_WRONG_COMPARTMENT (1468)
value ERROR_WRONG_DISK (34)
value ERROR_WRONG_EFS (6005)
value ERROR_WRONG_PASSWORD (1323)
value ERROR_WRONG_TARGET_NAME (1396)
value ERROR_XMLDSIG_ERROR (1466)
value ERROR_XML_ENCODING_MISMATCH (14100)
value ERROR_XML_PARSE_ERROR (1465)
value ESB_DISABLE_BOTH (0x0003)
value ESB_DISABLE_DOWN (0x0002)
value ESB_DISABLE_LEFT (0x0001)
value ESB_DISABLE_LTUP (ESB_DISABLE_LEFT)
value ESB_DISABLE_RIGHT (0x0002)
value ESB_DISABLE_RTDN (ESB_DISABLE_RIGHT)
value ESB_DISABLE_UP (0x0001)
value ESB_ENABLE_BOTH (0x0000)
value ESPIPE (29)
value ESRCH (3)
value ES_AUTOHSCROLL (0x0080L)
value ES_AUTOVSCROLL (0x0040L)
value ES_AWAYMODE_REQUIRED (((DWORD)0x00000040))
value ES_CENTER (0x0001L)
value ES_CONTINUOUS (((DWORD)0x80000000))
value ES_DISPLAY_REQUIRED (((DWORD)0x00000002))
value ES_LEFT (0x0000L)
value ES_LOWERCASE (0x0010L)
value ES_MULTILINE (0x0004L)
value ES_NOHIDESEL (0x0100L)
value ES_NUMBER (0x2000L)
value ES_OEMCONVERT (0x0400L)
value ES_PASSWORD (0x0020L)
value ES_READONLY (0x0800L)
value ES_RIGHT (0x0002L)
value ES_SYSTEM_REQUIRED (((DWORD)0x00000001))
value ES_UPPERCASE (0x0008L)
value ES_USER_PRESENT (((DWORD)0x00000004))
value ES_WANTRETURN (0x1000L)
value ETIME (137)
value ETIMEDOUT (138)
value ETO_CLIPPED (0x0004)
value ETO_GLYPH_INDEX (0x0010)
value ETO_IGNORELANGUAGE (0x1000)
value ETO_NUMERICSLATIN (0x0800)
value ETO_NUMERICSLOCAL (0x0400)
value ETO_OPAQUE (0x0002)
value ETO_PDY (0x2000)
value ETO_REVERSE_INDEX_MAP (0x10000)
value ETO_RTLREADING (0x0080)
value ETXTBSY (139)
value EVENPARITY (2)
value EVENTLOG_AUDIT_FAILURE (0x0010)
value EVENTLOG_AUDIT_SUCCESS (0x0008)
value EVENTLOG_BACKWARDS_READ (0x0008)
value EVENTLOG_END_ALL_PAIRED_EVENTS (0x0004)
value EVENTLOG_END_PAIRED_EVENT (0x0002)
value EVENTLOG_ERROR_TYPE (0x0001)
value EVENTLOG_FORWARDS_READ (0x0004)
value EVENTLOG_FULL_INFO (0)
value EVENTLOG_INFORMATION_TYPE (0x0004)
value EVENTLOG_PAIRED_EVENT_ACTIVE (0x0008)
value EVENTLOG_PAIRED_EVENT_INACTIVE (0x0010)
value EVENTLOG_SEEK_READ (0x0002)
value EVENTLOG_SEQUENTIAL_READ (0x0001)
value EVENTLOG_START_PAIRED_EVENT (0x0001)
value EVENTLOG_SUCCESS (0x0000)
value EVENTLOG_WARNING_TYPE (0x0002)
value EVENT_AIA_END (0xAFFF)
value EVENT_AIA_START (0xA000)
value EVENT_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED|SYNCHRONIZE|0x3))
value EVENT_CONSOLE_CARET (0x4001)
value EVENT_CONSOLE_END (0x40FF)
value EVENT_CONSOLE_END_APPLICATION (0x4007)
value EVENT_CONSOLE_LAYOUT (0x4005)
value EVENT_CONSOLE_START_APPLICATION (0x4006)
value EVENT_CONSOLE_UPDATE_REGION (0x4002)
value EVENT_CONSOLE_UPDATE_SCROLL (0x4004)
value EVENT_CONSOLE_UPDATE_SIMPLE (0x4003)
value EVENT_E_ALL_SUBSCRIBERS_FAILED (_HRESULT_TYPEDEF_(0x80040201L))
value EVENT_E_CANT_MODIFY_OR_DELETE_CONFIGURED_OBJECT (_HRESULT_TYPEDEF_(0x8004020EL))
value EVENT_E_CANT_MODIFY_OR_DELETE_UNCONFIGURED_OBJECT (_HRESULT_TYPEDEF_(0x8004020DL))
value EVENT_E_COMPLUS_NOT_INSTALLED (_HRESULT_TYPEDEF_(0x8004020CL))
value EVENT_E_FIRST (0x80040200L)
value EVENT_E_INTERNALERROR (_HRESULT_TYPEDEF_(0x80040206L))
value EVENT_E_INTERNALEXCEPTION (_HRESULT_TYPEDEF_(0x80040205L))
value EVENT_E_INVALID_EVENT_CLASS_PARTITION (_HRESULT_TYPEDEF_(0x8004020FL))
value EVENT_E_INVALID_PER_USER_SID (_HRESULT_TYPEDEF_(0x80040207L))
value EVENT_E_LAST (0x8004021FL)
value EVENT_E_MISSING_EVENTCLASS (_HRESULT_TYPEDEF_(0x8004020AL))
value EVENT_E_NOT_ALL_REMOVED (_HRESULT_TYPEDEF_(0x8004020BL))
value EVENT_E_PER_USER_SID_NOT_LOGGED_ON (_HRESULT_TYPEDEF_(0x80040210L))
value EVENT_E_QUERYFIELD (_HRESULT_TYPEDEF_(0x80040204L))
value EVENT_E_QUERYSYNTAX (_HRESULT_TYPEDEF_(0x80040203L))
value EVENT_E_TOO_MANY_METHODS (_HRESULT_TYPEDEF_(0x80040209L))
value EVENT_E_USER_EXCEPTION (_HRESULT_TYPEDEF_(0x80040208L))
value EVENT_MAX (0x7FFFFFFF)
value EVENT_MIN (0x00000001)
value EVENT_MODIFY_STATE (0x0002)
value EVENT_OBJECT_ACCELERATORCHANGE (0x8012)
value EVENT_OBJECT_CLOAKED (0x8017)
value EVENT_OBJECT_CONTENTSCROLLED (0x8015)
value EVENT_OBJECT_CREATE (0x8000)
value EVENT_OBJECT_DEFACTIONCHANGE (0x8011)
value EVENT_OBJECT_DESCRIPTIONCHANGE (0x800D)
value EVENT_OBJECT_DESTROY (0x8001)
value EVENT_OBJECT_DRAGCANCEL (0x8022)
value EVENT_OBJECT_DRAGCOMPLETE (0x8023)
value EVENT_OBJECT_DRAGDROPPED (0x8026)
value EVENT_OBJECT_DRAGENTER (0x8024)
value EVENT_OBJECT_DRAGLEAVE (0x8025)
value EVENT_OBJECT_DRAGSTART (0x8021)
value EVENT_OBJECT_END (0x80FF)
value EVENT_OBJECT_FOCUS (0x8005)
value EVENT_OBJECT_HELPCHANGE (0x8010)
value EVENT_OBJECT_HIDE (0x8003)
value EVENT_OBJECT_HOSTEDOBJECTSINVALIDATED (0x8020)
value EVENT_OBJECT_IME_CHANGE (0x8029)
value EVENT_OBJECT_IME_HIDE (0x8028)
value EVENT_OBJECT_IME_SHOW (0x8027)
value EVENT_OBJECT_INVOKED (0x8013)
value EVENT_OBJECT_LIVEREGIONCHANGED (0x8019)
value EVENT_OBJECT_LOCATIONCHANGE (0x800B)
value EVENT_OBJECT_NAMECHANGE (0x800C)
value EVENT_OBJECT_PARENTCHANGE (0x800F)
value EVENT_OBJECT_REORDER (0x8004)
value EVENT_OBJECT_SELECTION (0x8006)
value EVENT_OBJECT_SELECTIONADD (0x8007)
value EVENT_OBJECT_SELECTIONREMOVE (0x8008)
value EVENT_OBJECT_SELECTIONWITHIN (0x8009)
value EVENT_OBJECT_SHOW (0x8002)
value EVENT_OBJECT_STATECHANGE (0x800A)
value EVENT_OBJECT_TEXTEDIT_CONVERSIONTARGETCHANGED (0x8030)
value EVENT_OBJECT_TEXTSELECTIONCHANGED (0x8014)
value EVENT_OBJECT_UNCLOAKED (0x8018)
value EVENT_OBJECT_VALUECHANGE (0x800E)
value EVENT_OEM_DEFINED_END (0x01FF)
value EVENT_OEM_DEFINED_START (0x0101)
value EVENT_SYSTEM_ALERT (0x0002)
value EVENT_SYSTEM_ARRANGMENTPREVIEW (0x8016)
value EVENT_SYSTEM_CAPTUREEND (0x0009)
value EVENT_SYSTEM_CAPTURESTART (0x0008)
value EVENT_SYSTEM_CONTEXTHELPEND (0x000D)
value EVENT_SYSTEM_CONTEXTHELPSTART (0x000C)
value EVENT_SYSTEM_DESKTOPSWITCH (0x0020)
value EVENT_SYSTEM_DIALOGEND (0x0011)
value EVENT_SYSTEM_DIALOGSTART (0x0010)
value EVENT_SYSTEM_DRAGDROPEND (0x000F)
value EVENT_SYSTEM_DRAGDROPSTART (0x000E)
value EVENT_SYSTEM_END (0x00FF)
value EVENT_SYSTEM_FOREGROUND (0x0003)
value EVENT_SYSTEM_IME_KEY_NOTIFICATION (0x0029)
value EVENT_SYSTEM_MENUEND (0x0005)
value EVENT_SYSTEM_MENUPOPUPEND (0x0007)
value EVENT_SYSTEM_MENUPOPUPSTART (0x0006)
value EVENT_SYSTEM_MENUSTART (0x0004)
value EVENT_SYSTEM_MINIMIZEEND (0x0017)
value EVENT_SYSTEM_MINIMIZESTART (0x0016)
value EVENT_SYSTEM_MOVESIZEEND (0x000B)
value EVENT_SYSTEM_MOVESIZESTART (0x000A)
value EVENT_SYSTEM_SCROLLINGEND (0x0013)
value EVENT_SYSTEM_SCROLLINGSTART (0x0012)
value EVENT_SYSTEM_SOUND (0x0001)
value EVENT_SYSTEM_SWITCHEND (0x0015)
value EVENT_SYSTEM_SWITCHER_APPDROPPED (0x0026)
value EVENT_SYSTEM_SWITCHER_APPGRABBED (0x0024)
value EVENT_SYSTEM_SWITCHER_APPOVERTARGET (0x0025)
value EVENT_SYSTEM_SWITCHER_CANCELLED (0x0027)
value EVENT_SYSTEM_SWITCHSTART (0x0014)
value EVENT_S_FIRST (0x00040200L)
value EVENT_S_LAST (0x0004021FL)
value EVENT_S_NOSUBSCRIBERS (_HRESULT_TYPEDEF_(0x00040202L))
value EVENT_S_SOME_SUBSCRIBERS_FAILED (_HRESULT_TYPEDEF_(0x00040200L))
value EVENT_UIA_EVENTID_END (0x4EFF)
value EVENT_UIA_EVENTID_START (0x4E00)
value EVENT_UIA_PROPID_END (0x75FF)
value EVENT_UIA_PROPID_START (0x7500)
value EV_BREAK (0x0040)
value EV_CTS (0x0008)
value EV_DSR (0x0010)
value EV_ERR (0x0080)
value EV_PERR (0x0200)
value EV_RING (0x0100)
value EV_RLSD (0x0020)
value EV_RXCHAR (0x0001)
value EV_RXFLAG (0x0002)
value EV_TXEMPTY (0x0004)
value EWOULDBLOCK (140)
value EWX_ARSO (0x04000000)
value EWX_BOOTOPTIONS (0x01000000)
value EWX_CHECK_SAFE_FOR_SERVER (0x08000000)
value EWX_FORCE (0x00000004)
value EWX_FORCEIFHUNG (0x00000010)
value EWX_HYBRID_SHUTDOWN (0x00400000)
value EWX_LOGOFF (0x00000000)
value EWX_POWEROFF (0x00000008)
value EWX_QUICKRESOLVE (0x00000020)
value EWX_REBOOT (0x00000002)
value EWX_RESTARTAPPS (0x00000040)
value EWX_SHUTDOWN (0x00000001)
value EWX_SYSTEM_INITIATED (0x10000000)
value EXCEPTION_ACCESS_VIOLATION (STATUS_ACCESS_VIOLATION)
value EXCEPTION_ARRAY_BOUNDS_EXCEEDED (STATUS_ARRAY_BOUNDS_EXCEEDED)
value EXCEPTION_BREAKPOINT (STATUS_BREAKPOINT)
value EXCEPTION_COLLIDED_UNWIND (0x40)
value EXCEPTION_CONTINUE_EXECUTION ((-1))
value EXCEPTION_CONTINUE_SEARCH (0)
value EXCEPTION_DATATYPE_MISALIGNMENT (STATUS_DATATYPE_MISALIGNMENT)
value EXCEPTION_DEBUG_EVENT (1)
value EXCEPTION_EXECUTE_FAULT (8)
value EXCEPTION_EXECUTE_HANDLER (1)
value EXCEPTION_EXIT_UNWIND (0x4)
value EXCEPTION_FLT_DENORMAL_OPERAND (STATUS_FLOAT_DENORMAL_OPERAND)
value EXCEPTION_FLT_DIVIDE_BY_ZERO (STATUS_FLOAT_DIVIDE_BY_ZERO)
value EXCEPTION_FLT_INEXACT_RESULT (STATUS_FLOAT_INEXACT_RESULT)
value EXCEPTION_FLT_INVALID_OPERATION (STATUS_FLOAT_INVALID_OPERATION)
value EXCEPTION_FLT_OVERFLOW (STATUS_FLOAT_OVERFLOW)
value EXCEPTION_FLT_STACK_CHECK (STATUS_FLOAT_STACK_CHECK)
value EXCEPTION_FLT_UNDERFLOW (STATUS_FLOAT_UNDERFLOW)
value EXCEPTION_GUARD_PAGE (STATUS_GUARD_PAGE_VIOLATION)
value EXCEPTION_ILLEGAL_INSTRUCTION (STATUS_ILLEGAL_INSTRUCTION)
value EXCEPTION_INT_DIVIDE_BY_ZERO (STATUS_INTEGER_DIVIDE_BY_ZERO)
value EXCEPTION_INT_OVERFLOW (STATUS_INTEGER_OVERFLOW)
value EXCEPTION_INVALID_DISPOSITION (STATUS_INVALID_DISPOSITION)
value EXCEPTION_INVALID_HANDLE (STATUS_INVALID_HANDLE)
value EXCEPTION_IN_PAGE_ERROR (STATUS_IN_PAGE_ERROR)
value EXCEPTION_MAXIMUM_PARAMETERS (15)
value EXCEPTION_NESTED_CALL (0x10)
value EXCEPTION_NONCONTINUABLE (0x1)
value EXCEPTION_NONCONTINUABLE_EXCEPTION (STATUS_NONCONTINUABLE_EXCEPTION)
value EXCEPTION_POSSIBLE_DEADLOCK (STATUS_POSSIBLE_DEADLOCK)
value EXCEPTION_PRIV_INSTRUCTION (STATUS_PRIVILEGED_INSTRUCTION)
value EXCEPTION_READ_FAULT (0)
value EXCEPTION_SINGLE_STEP (STATUS_SINGLE_STEP)
value EXCEPTION_SOFTWARE_ORIGINATE (0x80)
value EXCEPTION_STACK_INVALID (0x8)
value EXCEPTION_STACK_OVERFLOW (STATUS_STACK_OVERFLOW)
value EXCEPTION_TARGET_UNWIND (0x20)
value EXCEPTION_UNWIND ((EXCEPTION_UNWINDING | EXCEPTION_EXIT_UNWIND | EXCEPTION_TARGET_UNWIND | EXCEPTION_COLLIDED_UNWIND))
value EXCEPTION_UNWINDING (0x2)
value EXCEPTION_WRITE_FAULT (1)
value EXDEV (18)
value EXECUTE_OFFLINE_DIAGS (0xD4)
value EXIT_FAILURE (1)
value EXIT_PROCESS_DEBUG_EVENT (5)
value EXIT_SUCCESS (0)
value EXIT_THREAD_DEBUG_EVENT (4)
value EXPENTRY (CALLBACK)
value EXPORT_PRIVATE_KEYS (0x0004)
value EXTENDED_STARTUPINFO_PRESENT (0x00080000)
value EXTEND_IEPORT (2)
value EXTTEXTOUT (512)
value EXT_DEVICE_CAPS (4099)
value E_ABORT (_HRESULT_TYPEDEF_(0x80004004L))
value E_ACCESSDENIED (_HRESULT_TYPEDEF_(0x80070005L))
value E_APPLICATION_ACTIVATION_EXEC_FAILURE (_HRESULT_TYPEDEF_(0x8027025BL))
value E_APPLICATION_ACTIVATION_TIMED_OUT (_HRESULT_TYPEDEF_(0x8027025AL))
value E_APPLICATION_EXITING (_HRESULT_TYPEDEF_(0x8000001AL))
value E_APPLICATION_MANAGER_NOT_RUNNING (_HRESULT_TYPEDEF_(0x80270257L))
value E_APPLICATION_NOT_REGISTERED (_HRESULT_TYPEDEF_(0x80270254L))
value E_APPLICATION_TEMPORARY_LICENSE_ERROR (_HRESULT_TYPEDEF_(0x8027025CL))
value E_APPLICATION_TRIAL_LICENSE_EXPIRED (_HRESULT_TYPEDEF_(0x8027025DL))
value E_APPLICATION_VIEW_EXITING (_HRESULT_TYPEDEF_(0x8000001BL))
value E_ASYNC_OPERATION_NOT_STARTED (_HRESULT_TYPEDEF_(0x80000019L))
value E_AUDIO_ENGINE_NODE_NOT_FOUND (_HRESULT_TYPEDEF_(0x80660001L))
value E_BLUETOOTH_ATT_ATTRIBUTE_NOT_FOUND (_HRESULT_TYPEDEF_(0x8065000AL))
value E_BLUETOOTH_ATT_ATTRIBUTE_NOT_LONG (_HRESULT_TYPEDEF_(0x8065000BL))
value E_BLUETOOTH_ATT_INSUFFICIENT_AUTHENTICATION (_HRESULT_TYPEDEF_(0x80650005L))
value E_BLUETOOTH_ATT_INSUFFICIENT_AUTHORIZATION (_HRESULT_TYPEDEF_(0x80650008L))
value E_BLUETOOTH_ATT_INSUFFICIENT_ENCRYPTION (_HRESULT_TYPEDEF_(0x8065000FL))
value E_BLUETOOTH_ATT_INSUFFICIENT_ENCRYPTION_KEY_SIZE (_HRESULT_TYPEDEF_(0x8065000CL))
value E_BLUETOOTH_ATT_INSUFFICIENT_RESOURCES (_HRESULT_TYPEDEF_(0x80650011L))
value E_BLUETOOTH_ATT_INVALID_ATTRIBUTE_VALUE_LENGTH (_HRESULT_TYPEDEF_(0x8065000DL))
value E_BLUETOOTH_ATT_INVALID_HANDLE (_HRESULT_TYPEDEF_(0x80650001L))
value E_BLUETOOTH_ATT_INVALID_OFFSET (_HRESULT_TYPEDEF_(0x80650007L))
value E_BLUETOOTH_ATT_INVALID_PDU (_HRESULT_TYPEDEF_(0x80650004L))
value E_BLUETOOTH_ATT_PREPARE_QUEUE_FULL (_HRESULT_TYPEDEF_(0x80650009L))
value E_BLUETOOTH_ATT_READ_NOT_PERMITTED (_HRESULT_TYPEDEF_(0x80650002L))
value E_BLUETOOTH_ATT_REQUEST_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80650006L))
value E_BLUETOOTH_ATT_UNKNOWN_ERROR (_HRESULT_TYPEDEF_(0x80651000L))
value E_BLUETOOTH_ATT_UNLIKELY (_HRESULT_TYPEDEF_(0x8065000EL))
value E_BLUETOOTH_ATT_UNSUPPORTED_GROUP_TYPE (_HRESULT_TYPEDEF_(0x80650010L))
value E_BLUETOOTH_ATT_WRITE_NOT_PERMITTED (_HRESULT_TYPEDEF_(0x80650003L))
value E_BOUNDS (_HRESULT_TYPEDEF_(0x8000000BL))
value E_CHANGED_STATE (_HRESULT_TYPEDEF_(0x8000000CL))
value E_DRAW (VIEW_E_DRAW)
value E_ELEVATED_ACTIVATION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80270251L))
value E_FAIL (_HRESULT_TYPEDEF_(0x80004005L))
value E_FULL_ADMIN_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80270253L))
value E_HANDLE (_HRESULT_TYPEDEF_(0x80070006L))
value E_HDAUDIO_CONNECTION_LIST_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80660003L))
value E_HDAUDIO_EMPTY_CONNECTION_LIST (_HRESULT_TYPEDEF_(0x80660002L))
value E_HDAUDIO_NO_LOGICAL_DEVICES_CREATED (_HRESULT_TYPEDEF_(0x80660004L))
value E_HDAUDIO_NULL_LINKED_LIST_ENTRY (_HRESULT_TYPEDEF_(0x80660005L))
value E_ILLEGAL_DELEGATE_ASSIGNMENT (_HRESULT_TYPEDEF_(0x80000018L))
value E_ILLEGAL_METHOD_CALL (_HRESULT_TYPEDEF_(0x8000000EL))
value E_ILLEGAL_STATE_CHANGE (_HRESULT_TYPEDEF_(0x8000000DL))
value E_INVALIDARG (_HRESULT_TYPEDEF_(0x80070057L))
value E_INVALID_PROTOCOL_FORMAT (_HRESULT_TYPEDEF_(0x83760002L))
value E_INVALID_PROTOCOL_OPERATION (_HRESULT_TYPEDEF_(0x83760001L))
value E_MBN_BAD_SIM (_HRESULT_TYPEDEF_(0x80548202L))
value E_MBN_CONTEXT_NOT_ACTIVATED (_HRESULT_TYPEDEF_(0x80548201L))
value E_MBN_DATA_CLASS_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x80548203L))
value E_MBN_DEFAULT_PROFILE_EXIST (_HRESULT_TYPEDEF_(0x80548219L))
value E_MBN_FAILURE (_HRESULT_TYPEDEF_(0x80548212L))
value E_MBN_INVALID_ACCESS_STRING (_HRESULT_TYPEDEF_(0x80548204L))
value E_MBN_INVALID_CACHE (_HRESULT_TYPEDEF_(0x8054820CL))
value E_MBN_INVALID_PROFILE (_HRESULT_TYPEDEF_(0x80548218L))
value E_MBN_MAX_ACTIVATED_CONTEXTS (_HRESULT_TYPEDEF_(0x80548205L))
value E_MBN_NOT_REGISTERED (_HRESULT_TYPEDEF_(0x8054820DL))
value E_MBN_PACKET_SVC_DETACHED (_HRESULT_TYPEDEF_(0x80548206L))
value E_MBN_PIN_DISABLED (_HRESULT_TYPEDEF_(0x80548211L))
value E_MBN_PIN_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8054820FL))
value E_MBN_PIN_REQUIRED (_HRESULT_TYPEDEF_(0x80548210L))
value E_MBN_PROVIDERS_NOT_FOUND (_HRESULT_TYPEDEF_(0x8054820EL))
value E_MBN_PROVIDER_NOT_VISIBLE (_HRESULT_TYPEDEF_(0x80548207L))
value E_MBN_RADIO_POWER_OFF (_HRESULT_TYPEDEF_(0x80548208L))
value E_MBN_SERVICE_NOT_ACTIVATED (_HRESULT_TYPEDEF_(0x80548209L))
value E_MBN_SIM_NOT_INSERTED (_HRESULT_TYPEDEF_(0x8054820AL))
value E_MBN_SMS_ENCODING_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80548220L))
value E_MBN_SMS_FILTER_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80548221L))
value E_MBN_SMS_FORMAT_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80548227L))
value E_MBN_SMS_INVALID_MEMORY_INDEX (_HRESULT_TYPEDEF_(0x80548222L))
value E_MBN_SMS_LANG_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80548223L))
value E_MBN_SMS_MEMORY_FAILURE (_HRESULT_TYPEDEF_(0x80548224L))
value E_MBN_SMS_MEMORY_FULL (_HRESULT_TYPEDEF_(0x80548229L))
value E_MBN_SMS_NETWORK_TIMEOUT (_HRESULT_TYPEDEF_(0x80548225L))
value E_MBN_SMS_OPERATION_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80548228L))
value E_MBN_SMS_UNKNOWN_SMSC_ADDRESS (_HRESULT_TYPEDEF_(0x80548226L))
value E_MBN_VOICE_CALL_IN_PROGRESS (_HRESULT_TYPEDEF_(0x8054820BL))
value E_MONITOR_RESOLUTION_TOO_LOW (_HRESULT_TYPEDEF_(0x80270250L))
value E_MULTIPLE_EXTENSIONS_FOR_APPLICATION (_HRESULT_TYPEDEF_(0x80270255L))
value E_MULTIPLE_PACKAGES_FOR_FAMILY (_HRESULT_TYPEDEF_(0x80270256L))
value E_NOINTERFACE (_HRESULT_TYPEDEF_(0x80004002L))
value E_NOTIMPL (_HRESULT_TYPEDEF_(0x80004001L))
value E_NOT_SET (HRESULT_FROM_WIN32(ERROR_NOT_FOUND))
value E_NOT_SUFFICIENT_BUFFER (HRESULT_FROM_WIN32(ERROR_INSUFFICIENT_BUFFER))
value E_NOT_VALID_STATE (HRESULT_FROM_WIN32(ERROR_INVALID_STATE))
value E_NO_TASK_QUEUE (HRESULT_FROM_WIN32(ERROR_NO_TASK_QUEUE))
value E_OUTOFMEMORY (_HRESULT_TYPEDEF_(0x8007000EL))
value E_PENDING (_HRESULT_TYPEDEF_(0x8000000AL))
value E_POINTER (_HRESULT_TYPEDEF_(0x80004003L))
value E_PROTOCOL_EXTENSIONS_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x83760003L))
value E_PROTOCOL_VERSION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x83760005L))
value E_SKYDRIVE_FILE_NOT_UPLOADED (_HRESULT_TYPEDEF_(0x80270263L))
value E_SKYDRIVE_ROOT_TARGET_CANNOT_INDEX (_HRESULT_TYPEDEF_(0x80270262L))
value E_SKYDRIVE_ROOT_TARGET_FILE_SYSTEM_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80270260L))
value E_SKYDRIVE_ROOT_TARGET_OVERLAP (_HRESULT_TYPEDEF_(0x80270261L))
value E_SKYDRIVE_ROOT_TARGET_VOLUME_ROOT_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80270265L))
value E_SKYDRIVE_UPDATE_AVAILABILITY_FAIL (_HRESULT_TYPEDEF_(0x80270264L))
value E_STRING_NOT_NULL_TERMINATED (_HRESULT_TYPEDEF_(0x80000017L))
value E_SUBPROTOCOL_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x83760004L))
value E_SYNCENGINE_CLIENT_UPDATE_NEEDED (_HRESULT_TYPEDEF_(0x8802D006L))
value E_SYNCENGINE_FILE_IDENTIFIER_UNKNOWN (_HRESULT_TYPEDEF_(0x8802C002L))
value E_SYNCENGINE_FILE_SIZE_EXCEEDS_REMAINING_QUOTA (_HRESULT_TYPEDEF_(0x8802B002L))
value E_SYNCENGINE_FILE_SIZE_OVER_LIMIT (_HRESULT_TYPEDEF_(0x8802B001L))
value E_SYNCENGINE_FILE_SYNC_PARTNER_ERROR (_HRESULT_TYPEDEF_(0x8802B005L))
value E_SYNCENGINE_FOLDER_INACCESSIBLE (_HRESULT_TYPEDEF_(0x8802D001L))
value E_SYNCENGINE_FOLDER_IN_REDIRECTION (_HRESULT_TYPEDEF_(0x8802D00BL))
value E_SYNCENGINE_FOLDER_ITEM_COUNT_LIMIT_EXCEEDED (_HRESULT_TYPEDEF_(0x8802B004L))
value E_SYNCENGINE_PATH_LENGTH_LIMIT_EXCEEDED (_HRESULT_TYPEDEF_(0x8802D004L))
value E_SYNCENGINE_PROXY_AUTHENTICATION_REQUIRED (_HRESULT_TYPEDEF_(0x8802D007L))
value E_SYNCENGINE_REMOTE_PATH_LENGTH_LIMIT_EXCEEDED (_HRESULT_TYPEDEF_(0x8802D005L))
value E_SYNCENGINE_REQUEST_BLOCKED_BY_SERVICE (_HRESULT_TYPEDEF_(0x8802C006L))
value E_SYNCENGINE_REQUEST_BLOCKED_DUE_TO_CLIENT_ERROR (_HRESULT_TYPEDEF_(0x8802C007L))
value E_SYNCENGINE_SERVICE_AUTHENTICATION_FAILED (_HRESULT_TYPEDEF_(0x8802C003L))
value E_SYNCENGINE_SERVICE_RETURNED_UNEXPECTED_SIZE (_HRESULT_TYPEDEF_(0x8802C005L))
value E_SYNCENGINE_STORAGE_SERVICE_BLOCKED (_HRESULT_TYPEDEF_(0x8802D00AL))
value E_SYNCENGINE_STORAGE_SERVICE_PROVISIONING_FAILED (_HRESULT_TYPEDEF_(0x8802D008L))
value E_SYNCENGINE_SYNC_PAUSED_BY_SERVICE (_HRESULT_TYPEDEF_(0x8802B006L))
value E_SYNCENGINE_UNKNOWN_SERVICE_ERROR (_HRESULT_TYPEDEF_(0x8802C004L))
value E_SYNCENGINE_UNSUPPORTED_FILE_NAME (_HRESULT_TYPEDEF_(0x8802B003L))
value E_SYNCENGINE_UNSUPPORTED_FOLDER_NAME (_HRESULT_TYPEDEF_(0x8802D002L))
value E_SYNCENGINE_UNSUPPORTED_MARKET (_HRESULT_TYPEDEF_(0x8802D003L))
value E_SYNCENGINE_UNSUPPORTED_REPARSE_POINT (_HRESULT_TYPEDEF_(0x8802D009L))
value E_TIME_SENSITIVE_THREAD (HRESULT_FROM_WIN32(ERROR_TIME_SENSITIVE_THREAD))
value E_UAC_DISABLED (_HRESULT_TYPEDEF_(0x80270252L))
value E_UNEXPECTED (_HRESULT_TYPEDEF_(0x8000FFFFL))
value FACILITY_AAF (18)
value FACILITY_ACCELERATOR (1536)
value FACILITY_ACS (20)
value FACILITY_ACTION_QUEUE (44)
value FACILITY_AUDCLNT (2185)
value FACILITY_AUDIO (102)
value FACILITY_AUDIOSTREAMING (1094)
value FACILITY_BACKGROUNDCOPY (32)
value FACILITY_BCD (57)
value FACILITY_BLB (120)
value FACILITY_BLBUI (128)
value FACILITY_BLB_CLI (121)
value FACILITY_BLUETOOTH_ATT (101)
value FACILITY_CERT (11)
value FACILITY_CMI (54)
value FACILITY_COMPLUS (17)
value FACILITY_CONFIGURATION (33)
value FACILITY_CONTROL (10)
value FACILITY_DAF (100)
value FACILITY_DEBUGGERS (176)
value FACILITY_DEFRAG (2304)
value FACILITY_DELIVERY_OPTIMIZATION (208)
value FACILITY_DEPLOYMENT_SERVICES_BINLSVC (261)
value FACILITY_DEPLOYMENT_SERVICES_CONTENT_PROVIDER (293)
value FACILITY_DEPLOYMENT_SERVICES_DRIVER_PROVISIONING (278)
value FACILITY_DEPLOYMENT_SERVICES_IMAGING (258)
value FACILITY_DEPLOYMENT_SERVICES_MANAGEMENT (259)
value FACILITY_DEPLOYMENT_SERVICES_MULTICAST_CLIENT (290)
value FACILITY_DEPLOYMENT_SERVICES_MULTICAST_SERVER (289)
value FACILITY_DEPLOYMENT_SERVICES_PXE (263)
value FACILITY_DEPLOYMENT_SERVICES_SERVER (257)
value FACILITY_DEPLOYMENT_SERVICES_TFTP (264)
value FACILITY_DEPLOYMENT_SERVICES_TRANSPORT_MANAGEMENT (272)
value FACILITY_DEPLOYMENT_SERVICES_UTIL (260)
value FACILITY_DEVICE_UPDATE_AGENT (135)
value FACILITY_DIRECTMUSIC (2168)
value FACILITY_DIRECTORYSERVICE (37)
value FACILITY_DISPATCH (2)
value FACILITY_DLS (153)
value FACILITY_DMSERVER (256)
value FACILITY_DPLAY (21)
value FACILITY_DRVSERVICING (136)
value FACILITY_DXCORE (2176)
value FACILITY_DXGI (2170)
value FACILITY_DXGI_DDI (2171)
value FACILITY_EAP (66)
value FACILITY_EAS (85)
value FACILITY_FVE (49)
value FACILITY_FWP (50)
value FACILITY_GAME (2340)
value FACILITY_GRAPHICS (38)
value FACILITY_HSP_SERVICES (296)
value FACILITY_HSP_SOFTWARE (297)
value FACILITY_HTTP (25)
value FACILITY_INPUT (64)
value FACILITY_INTERNET (12)
value FACILITY_IORING (70)
value FACILITY_ITF (4)
value FACILITY_JSCRIPT (2306)
value FACILITY_LEAP (2184)
value FACILITY_LINGUISTIC_SERVICES (305)
value FACILITY_MBN (84)
value FACILITY_MEDIASERVER (13)
value FACILITY_METADIRECTORY (35)
value FACILITY_MOBILE (1793)
value FACILITY_MSMQ (14)
value FACILITY_NAP (39)
value FACILITY_NDIS (52)
value FACILITY_NT_BIT (0x10000000)
value FACILITY_NULL (0)
value FACILITY_OCP_UPDATE_AGENT (173)
value FACILITY_ONLINE_ID (134)
value FACILITY_OPC (81)
value FACILITY_PARSE (113)
value FACILITY_PIDGENX (2561)
value FACILITY_PIX (2748)
value FACILITY_PLA (48)
value FACILITY_POWERSHELL (84)
value FACILITY_PRESENTATION (2177)
value FACILITY_QUIC (65)
value FACILITY_RAS (83)
value FACILITY_RESTORE (256)
value FACILITY_RPC (1)
value FACILITY_SCARD (16)
value FACILITY_SCRIPT (112)
value FACILITY_SDIAG (60)
value FACILITY_SECURITY (9)
value FACILITY_SERVICE_FABRIC (1968)
value FACILITY_SETUPAPI (15)
value FACILITY_SHELL (39)
value FACILITY_SOS (160)
value FACILITY_SPP (256)
value FACILITY_SQLITE (1967)
value FACILITY_SSPI (9)
value FACILITY_STATEREPOSITORY (103)
value FACILITY_STATE_MANAGEMENT (34)
value FACILITY_STORAGE (3)
value FACILITY_SXS (23)
value FACILITY_SYNCENGINE (2050)
value FACILITY_TIERING (131)
value FACILITY_TPM_SERVICES (40)
value FACILITY_TPM_SOFTWARE (41)
value FACILITY_TTD (1490)
value FACILITY_UI (42)
value FACILITY_UMI (22)
value FACILITY_URT (19)
value FACILITY_USERMODE_COMMONLOG (26)
value FACILITY_USERMODE_FILTER_MANAGER (31)
value FACILITY_USERMODE_HNS (59)
value FACILITY_USERMODE_HYPERVISOR (53)
value FACILITY_USERMODE_LICENSING (234)
value FACILITY_USERMODE_SDBUS (2305)
value FACILITY_USERMODE_SPACES (231)
value FACILITY_USERMODE_VHD (58)
value FACILITY_USERMODE_VIRTUALIZATION (55)
value FACILITY_USERMODE_VOLMGR (56)
value FACILITY_USERMODE_VOLSNAP (130)
value FACILITY_USER_MODE_SECURITY_CORE (232)
value FACILITY_USN (129)
value FACILITY_UTC (1989)
value FACILITY_VISUALCPP (109)
value FACILITY_WEB (885)
value FACILITY_WEBSERVICES (61)
value FACILITY_WEB_SOCKET (886)
value FACILITY_WEP (2049)
value FACILITY_WER (27)
value FACILITY_WIA (33)
value FACILITY_WINCODEC_DWRITE_DWM (2200)
value FACILITY_WINDOWS (8)
value FACILITY_WINDOWSUPDATE (36)
value FACILITY_WINDOWS_CE (24)
value FACILITY_WINDOWS_DEFENDER (80)
value FACILITY_WINDOWS_SETUP (48)
value FACILITY_WINDOWS_STORE (63)
value FACILITY_WINML (2192)
value FACILITY_WINPE (61)
value FACILITY_WINRM (51)
value FACILITY_WMAAECMA (1996)
value FACILITY_WPN (62)
value FACILITY_WSBAPP (122)
value FACILITY_WSB_ONLINE (133)
value FACILITY_XAML (43)
value FACILITY_XBOX (2339)
value FACILITY_XPS (82)
value FADF_AUTO (( 0x1 ))
value FADF_BSTR (( 0x100 ))
value FADF_DISPATCH (( 0x400 ))
value FADF_EMBEDDED (( 0x4 ))
value FADF_FIXEDSIZE (( 0x10 ))
value FADF_HAVEIID (( 0x40 ))
value FADF_HAVEVARTYPE (( 0x80 ))
value FADF_RECORD (( 0x20 ))
value FADF_STATIC (( 0x2 ))
value FADF_UNKNOWN (( 0x200 ))
value FADF_VARIANT (( 0x800 ))
value FAILED_ACCESS_ACE_FLAG ((0x80))
value FAIL_FAST_GENERATE_EXCEPTION_ADDRESS (0x1)
value FAIL_FAST_NO_HARD_ERROR_DLG (0x2)
value FALSE (0)
value FALT (0x10)
value FAPPCOMMAND_KEY (0)
value FAPPCOMMAND_MASK (0xF000)
value FAPPCOMMAND_MOUSE (0x8000)
value FAPPCOMMAND_OEM (0x1000)
value FAST_FAIL_ADMINLESS_ACCESS_DENIED (55)
value FAST_FAIL_APCS_DISABLED (32)
value FAST_FAIL_CAST_GUARD (65)
value FAST_FAIL_CERTIFICATION_FAILURE (20)
value FAST_FAIL_CONTROL_INVALID_RETURN_ADDRESS (57)
value FAST_FAIL_CORRUPT_LIST_ENTRY (3)
value FAST_FAIL_CRYPTO_LIBRARY (22)
value FAST_FAIL_DEPRECATED_SERVICE_INVOKED (27)
value FAST_FAIL_DLOAD_PROTECTION_FAILURE (25)
value FAST_FAIL_ENCLAVE_CALL_FAILURE (53)
value FAST_FAIL_ETW_CORRUPTION (61)
value FAST_FAIL_FATAL_APP_EXIT (7)
value FAST_FAIL_FLAGS_CORRUPTION (59)
value FAST_FAIL_GS_COOKIE_INIT (6)
value FAST_FAIL_GUARD_EXPORT_SUPPRESSION_FAILURE (46)
value FAST_FAIL_GUARD_ICALL_CHECK_FAILURE (10)
value FAST_FAIL_GUARD_ICALL_CHECK_FAILURE_XFG (64)
value FAST_FAIL_GUARD_ICALL_CHECK_SUPPRESSED (31)
value FAST_FAIL_GUARD_JUMPTABLE (37)
value FAST_FAIL_GUARD_SS_FAILURE (44)
value FAST_FAIL_GUARD_WRITE_CHECK_FAILURE (11)
value FAST_FAIL_HEAP_METADATA_CORRUPTION (50)
value FAST_FAIL_HOST_VISIBILITY_CHANGE (66)
value FAST_FAIL_INCORRECT_STACK (4)
value FAST_FAIL_INVALID_ARG (5)
value FAST_FAIL_INVALID_BALANCED_TREE (29)
value FAST_FAIL_INVALID_BUFFER_ACCESS (28)
value FAST_FAIL_INVALID_CALL_IN_DLL_CALLOUT (23)
value FAST_FAIL_INVALID_CONTROL_STACK (47)
value FAST_FAIL_INVALID_DISPATCH_CONTEXT (39)
value FAST_FAIL_INVALID_EXCEPTION_CHAIN (21)
value FAST_FAIL_INVALID_FAST_FAIL_CODE (0xFFFFFFFF)
value FAST_FAIL_INVALID_FIBER_SWITCH (12)
value FAST_FAIL_INVALID_FILE_OPERATION (42)
value FAST_FAIL_INVALID_FLS_DATA (70)
value FAST_FAIL_INVALID_IAT (49)
value FAST_FAIL_INVALID_IDLE_STATE (33)
value FAST_FAIL_INVALID_IMAGE_BASE (24)
value FAST_FAIL_INVALID_JUMP_BUFFER (18)
value FAST_FAIL_INVALID_LOCK_STATE (36)
value FAST_FAIL_INVALID_LONGJUMP_TARGET (38)
value FAST_FAIL_INVALID_NEXT_THREAD (30)
value FAST_FAIL_INVALID_PFN (63)
value FAST_FAIL_INVALID_REFERENCE_COUNT (14)
value FAST_FAIL_INVALID_SET_OF_CONTEXT (13)
value FAST_FAIL_INVALID_SYSCALL_NUMBER (41)
value FAST_FAIL_INVALID_THREAD (40)
value FAST_FAIL_KERNEL_CET_SHADOW_STACK_ASSIST (67)
value FAST_FAIL_LEGACY_GS_VIOLATION (0)
value FAST_FAIL_LOADER_CONTINUITY_FAILURE (45)
value FAST_FAIL_LOW_LABEL_ACCESS_DENIED (52)
value FAST_FAIL_LPAC_ACCESS_DENIED (43)
value FAST_FAIL_MRDATA_MODIFIED (19)
value FAST_FAIL_MRDATA_PROTECTION_FAILURE (34)
value FAST_FAIL_NTDLL_PATCH_FAILED (69)
value FAST_FAIL_PATCH_CALLBACK_FAILED (68)
value FAST_FAIL_PAYLOAD_RESTRICTION_VIOLATION (51)
value FAST_FAIL_RANGE_CHECK_FAILURE (8)
value FAST_FAIL_RIO_ABORT (62)
value FAST_FAIL_SET_CONTEXT_DENIED (48)
value FAST_FAIL_STACK_COOKIE_CHECK_FAILURE (2)
value FAST_FAIL_UNEXPECTED_CALL (56)
value FAST_FAIL_UNEXPECTED_HEAP_EXCEPTION (35)
value FAST_FAIL_UNEXPECTED_HOST_BEHAVIOR (58)
value FAST_FAIL_UNHANDLED_LSS_EXCEPTON (54)
value FAST_FAIL_UNSAFE_EXTENSION_CALL (26)
value FAST_FAIL_UNSAFE_REGISTRY_ACCESS (9)
value FAST_FAIL_VEH_CORRUPTION (60)
value FAST_FAIL_VTGUARD_CHECK_FAILURE (1)
value FA_E_HOMEGROUP_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x80270222L))
value FA_E_MAX_PERSISTED_ITEMS_REACHED (_HRESULT_TYPEDEF_(0x80270220L))
value FCONTROL (0x08)
value FD_ACCEPT_BIT (3)
value FD_ADDRESS_LIST_CHANGE_BIT (9)
value FD_CLOSE_BIT (5)
value FD_CONNECT_BIT (4)
value FD_GROUP_QOS_BIT (7)
value FD_MAX_EVENTS (10)
value FD_OOB_BIT (2)
value FD_QOS_BIT (6)
value FD_READ_BIT (0)
value FD_ROUTING_INTERFACE_CHANGE_BIT (8)
value FD_SETSIZE (64)
value FD_WRITE_BIT (1)
value FEATURESETTING_CUSTPAPER (3)
value FEATURESETTING_MIRROR (4)
value FEATURESETTING_NEGATIVE (5)
value FEATURESETTING_NUP (0)
value FEATURESETTING_OUTPUT (1)
value FEATURESETTING_PRIVATE_BEGIN (0x1000)
value FEATURESETTING_PRIVATE_END (0x1FFF)
value FEATURESETTING_PROTOCOL (6)
value FEATURESETTING_PSLEVEL (2)
value FE_FONTSMOOTHINGCLEARTYPE (0x0002)
value FE_FONTSMOOTHINGORIENTATIONBGR (0x0000)
value FE_FONTSMOOTHINGORIENTATIONRGB (0x0001)
value FE_FONTSMOOTHINGSTANDARD (0x0001)
value FIBER_FLAG_FLOAT_SWITCH (0x1)
value FIEF_FLAG_FORCE_JITUI (0x1)
value FIEF_FLAG_PEEK (0x2)
value FIEF_FLAG_SKIP_INSTALLED_VERSION_CHECK (0x4)
value FILENAME_MAX (260)
value FILEOKSTRING (FILEOKSTRINGA)
value FILEOPENORD (1536)
value FILESYSTEM_STATISTICS_TYPE_EXFAT (3)
value FILESYSTEM_STATISTICS_TYPE_FAT (2)
value FILESYSTEM_STATISTICS_TYPE_NTFS (1)
value FILESYSTEM_STATISTICS_TYPE_REFS (4)
value FILE_ACTION_ADDED (0x00000001)
value FILE_ACTION_MODIFIED (0x00000003)
value FILE_ACTION_REMOVED (0x00000002)
value FILE_ACTION_RENAMED_NEW_NAME (0x00000005)
value FILE_ACTION_RENAMED_OLD_NAME (0x00000004)
value FILE_ADD_FILE (( 0x0002 ))
value FILE_ADD_SUBDIRECTORY (( 0x0004 ))
value FILE_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | SYNCHRONIZE | 0x1FF))
value FILE_ANY_ACCESS (0)
value FILE_APPEND_DATA (( 0x0004 ))
value FILE_ATTRIBUTE_ARCHIVE (0x00000020)
value FILE_ATTRIBUTE_COMPRESSED (0x00000800)
value FILE_ATTRIBUTE_DEVICE (0x00000040)
value FILE_ATTRIBUTE_DIRECTORY (0x00000010)
value FILE_ATTRIBUTE_EA (0x00040000)
value FILE_ATTRIBUTE_ENCRYPTED (0x00004000)
value FILE_ATTRIBUTE_HIDDEN (0x00000002)
value FILE_ATTRIBUTE_INTEGRITY_STREAM (0x00008000)
value FILE_ATTRIBUTE_NORMAL (0x00000080)
value FILE_ATTRIBUTE_NOT_CONTENT_INDEXED (0x00002000)
value FILE_ATTRIBUTE_NO_SCRUB_DATA (0x00020000)
value FILE_ATTRIBUTE_OFFLINE (0x00001000)
value FILE_ATTRIBUTE_PINNED (0x00080000)
value FILE_ATTRIBUTE_READONLY (0x00000001)
value FILE_ATTRIBUTE_RECALL_ON_DATA_ACCESS (0x00400000)
value FILE_ATTRIBUTE_RECALL_ON_OPEN (0x00040000)
value FILE_ATTRIBUTE_REPARSE_POINT (0x00000400)
value FILE_ATTRIBUTE_SPARSE_FILE (0x00000200)
value FILE_ATTRIBUTE_STRICTLY_SEQUENTIAL (0x20000000)
value FILE_ATTRIBUTE_SYSTEM (0x00000004)
value FILE_ATTRIBUTE_TEMPORARY (0x00000100)
value FILE_ATTRIBUTE_UNPINNED (0x00100000)
value FILE_ATTRIBUTE_VIRTUAL (0x00010000)
value FILE_BEGIN (0)
value FILE_CACHE_MAX_HARD_DISABLE (0x00000002)
value FILE_CACHE_MAX_HARD_ENABLE (0x00000001)
value FILE_CACHE_MIN_HARD_DISABLE (0x00000008)
value FILE_CACHE_MIN_HARD_ENABLE (0x00000004)
value FILE_CASE_PRESERVED_NAMES (0x00000002)
value FILE_CASE_SENSITIVE_SEARCH (0x00000001)
value FILE_CLEAR_ENCRYPTION (0x00000002)
value FILE_CREATE_PIPE_INSTANCE (( 0x0004 ))
value FILE_CS_FLAG_CASE_SENSITIVE_DIR (0x00000001)
value FILE_CURRENT (1)
value FILE_DAX_VOLUME (0x20000000)
value FILE_DELETE_CHILD (( 0x0040 ))
value FILE_DEVICE_ACPI (0x00000032)
value FILE_DEVICE_BATTERY (0x00000029)
value FILE_DEVICE_BEEP (0x00000001)
value FILE_DEVICE_BIOMETRIC (0x00000044)
value FILE_DEVICE_BLUETOOTH (0x00000041)
value FILE_DEVICE_BUS_EXTENDER (0x0000002a)
value FILE_DEVICE_CD_ROM (0x00000002)
value FILE_DEVICE_CD_ROM_FILE_SYSTEM (0x00000003)
value FILE_DEVICE_CHANGER (0x00000030)
value FILE_DEVICE_CONSOLE (0x00000050)
value FILE_DEVICE_CONTROLLER (0x00000004)
value FILE_DEVICE_CRYPT_PROVIDER (0x0000003F)
value FILE_DEVICE_DATALINK (0x00000005)
value FILE_DEVICE_DEVAPI (0x00000047)
value FILE_DEVICE_DFS (0x00000006)
value FILE_DEVICE_DFS_FILE_SYSTEM (0x00000035)
value FILE_DEVICE_DFS_VOLUME (0x00000036)
value FILE_DEVICE_DISK (0x00000007)
value FILE_DEVICE_DISK_FILE_SYSTEM (0x00000008)
value FILE_DEVICE_DVD (0x00000033)
value FILE_DEVICE_EHSTOR (0x00000046)
value FILE_DEVICE_EVENT_COLLECTOR (0x0000005f)
value FILE_DEVICE_FILE_SYSTEM (0x00000009)
value FILE_DEVICE_FIPS (0x0000003A)
value FILE_DEVICE_FULLSCREEN_VIDEO (0x00000034)
value FILE_DEVICE_GPIO (0x00000048)
value FILE_DEVICE_HOLOGRAPHIC (0x0000005b)
value FILE_DEVICE_INFINIBAND (0x0000003B)
value FILE_DEVICE_INPORT_PORT (0x0000000a)
value FILE_DEVICE_KEYBOARD (0x0000000b)
value FILE_DEVICE_KS (0x0000002f)
value FILE_DEVICE_KSEC (0x00000039)
value FILE_DEVICE_MAILSLOT (0x0000000c)
value FILE_DEVICE_MASS_STORAGE (0x0000002d)
value FILE_DEVICE_MIDI_IN (0x0000000d)
value FILE_DEVICE_MIDI_OUT (0x0000000e)
value FILE_DEVICE_MODEM (0x0000002b)
value FILE_DEVICE_MOUSE (0x0000000f)
value FILE_DEVICE_MT_COMPOSITE (0x00000042)
value FILE_DEVICE_MT_TRANSPORT (0x00000043)
value FILE_DEVICE_MULTI_UNC_PROVIDER (0x00000010)
value FILE_DEVICE_NAMED_PIPE (0x00000011)
value FILE_DEVICE_NETWORK (0x00000012)
value FILE_DEVICE_NETWORK_BROWSER (0x00000013)
value FILE_DEVICE_NETWORK_FILE_SYSTEM (0x00000014)
value FILE_DEVICE_NETWORK_REDIRECTOR (0x00000028)
value FILE_DEVICE_NFP (0x00000051)
value FILE_DEVICE_NULL (0x00000015)
value FILE_DEVICE_NVDIMM (0x0000005a)
value FILE_DEVICE_PARALLEL_PORT (0x00000016)
value FILE_DEVICE_PERSISTENT_MEMORY (0x00000059)
value FILE_DEVICE_PHYSICAL_NETCARD (0x00000017)
value FILE_DEVICE_PMI (0x00000045)
value FILE_DEVICE_POINT_OF_SERVICE (0x00000054)
value FILE_DEVICE_PRINTER (0x00000018)
value FILE_DEVICE_PRM (0x0000005e)
value FILE_DEVICE_SCANNER (0x00000019)
value FILE_DEVICE_SCREEN (0x0000001c)
value FILE_DEVICE_SDFXHCI (0x0000005c)
value FILE_DEVICE_SERENUM (0x00000037)
value FILE_DEVICE_SERIAL_MOUSE_PORT (0x0000001a)
value FILE_DEVICE_SERIAL_PORT (0x0000001b)
value FILE_DEVICE_SMARTCARD (0x00000031)
value FILE_DEVICE_SMB (0x0000002e)
value FILE_DEVICE_SOUND (0x0000001d)
value FILE_DEVICE_SOUNDWIRE (0x00000061)
value FILE_DEVICE_STORAGE_REPLICATION (0x00000055)
value FILE_DEVICE_STREAMS (0x0000001e)
value FILE_DEVICE_SYSENV (0x00000052)
value FILE_DEVICE_TAPE (0x0000001f)
value FILE_DEVICE_TAPE_FILE_SYSTEM (0x00000020)
value FILE_DEVICE_TERMSRV (0x00000038)
value FILE_DEVICE_TRANSPORT (0x00000021)
value FILE_DEVICE_TRUST_ENV (0x00000056)
value FILE_DEVICE_UCM (0x00000057)
value FILE_DEVICE_UCMTCPCI (0x00000058)
value FILE_DEVICE_UCMUCSI (0x0000005d)
value FILE_DEVICE_UNKNOWN (0x00000022)
value FILE_DEVICE_USBEX (0x00000049)
value FILE_DEVICE_VDM (0x0000002c)
value FILE_DEVICE_VIDEO (0x00000023)
value FILE_DEVICE_VIRTUAL_BLOCK (0x00000053)
value FILE_DEVICE_VIRTUAL_DISK (0x00000024)
value FILE_DEVICE_VMBUS (0x0000003E)
value FILE_DEVICE_WAVE_IN (0x00000025)
value FILE_DEVICE_WAVE_OUT (0x00000026)
value FILE_DEVICE_WPD (0x00000040)
value FILE_DIR_DISALLOWED (9)
value FILE_DISPOSITION_FLAG_DELETE (0x00000001)
value FILE_DISPOSITION_FLAG_DO_NOT_DELETE (0x00000000)
value FILE_DISPOSITION_FLAG_FORCE_IMAGE_SECTION_CHECK (0x00000004)
value FILE_DISPOSITION_FLAG_IGNORE_READONLY_ATTRIBUTE (0x00000010)
value FILE_DISPOSITION_FLAG_ON_CLOSE (0x00000008)
value FILE_DISPOSITION_FLAG_POSIX_SEMANTICS (0x00000002)
value FILE_ENCRYPTABLE (0)
value FILE_END (2)
value FILE_EXECUTE (( 0x0020 ))
value FILE_FILE_COMPRESSION (0x00000010)
value FILE_FLAG_BACKUP_SEMANTICS (0x02000000)
value FILE_FLAG_DELETE_ON_CLOSE (0x04000000)
value FILE_FLAG_FIRST_PIPE_INSTANCE (0x00080000)
value FILE_FLAG_NO_BUFFERING (0x20000000)
value FILE_FLAG_OPEN_NO_RECALL (0x00100000)
value FILE_FLAG_OPEN_REPARSE_POINT (0x00200000)
value FILE_FLAG_OPEN_REQUIRING_OPLOCK (0x00040000)
value FILE_FLAG_OVERLAPPED (0x40000000)
value FILE_FLAG_POSIX_SEMANTICS (0x01000000)
value FILE_FLAG_RANDOM_ACCESS (0x10000000)
value FILE_FLAG_SEQUENTIAL_SCAN (0x08000000)
value FILE_FLAG_SESSION_AWARE (0x00800000)
value FILE_FLAG_WRITE_THROUGH (0x80000000)
value FILE_GENERIC_EXECUTE ((STANDARD_RIGHTS_EXECUTE | FILE_READ_ATTRIBUTES | FILE_EXECUTE | SYNCHRONIZE))
value FILE_GENERIC_READ ((STANDARD_RIGHTS_READ | FILE_READ_DATA | FILE_READ_ATTRIBUTES | FILE_READ_EA | SYNCHRONIZE))
value FILE_GENERIC_WRITE ((STANDARD_RIGHTS_WRITE | FILE_WRITE_DATA | FILE_WRITE_ATTRIBUTES | FILE_WRITE_EA | FILE_APPEND_DATA | SYNCHRONIZE))
value FILE_INVALID_FILE_ID (((LONGLONG)-1LL))
value FILE_IS_ENCRYPTED (1)
value FILE_LAYOUT_NAME_ENTRY_DOS ((0x00000002))
value FILE_LAYOUT_NAME_ENTRY_PRIMARY ((0x00000001))
value FILE_LIST_DIRECTORY (( 0x0001 ))
value FILE_MAP_ALL_ACCESS (SECTION_ALL_ACCESS)
value FILE_MAP_COPY (0x00000001)
value FILE_MAP_EXECUTE (SECTION_MAP_EXECUTE_EXPLICIT)
value FILE_MAP_LARGE_PAGES (0x20000000)
value FILE_MAP_READ (SECTION_MAP_READ)
value FILE_MAP_RESERVE (0x80000000)
value FILE_MAP_TARGETS_INVALID (0x40000000)
value FILE_MAP_WRITE (SECTION_MAP_WRITE)
value FILE_NAMED_STREAMS (0x00040000)
value FILE_NAME_FLAGS_UNSPECIFIED (0x80)
value FILE_NAME_FLAG_BOTH (0x03)
value FILE_NAME_FLAG_DOS (0x02)
value FILE_NAME_FLAG_HARDLINK (0)
value FILE_NAME_FLAG_NTFS (0x01)
value FILE_NAME_NORMALIZED (0x0)
value FILE_NAME_OPENED (0x8)
value FILE_NOTIFY_CHANGE_ATTRIBUTES (0x00000004)
value FILE_NOTIFY_CHANGE_CREATION (0x00000040)
value FILE_NOTIFY_CHANGE_DIR_NAME (0x00000002)
value FILE_NOTIFY_CHANGE_FILE_NAME (0x00000001)
value FILE_NOTIFY_CHANGE_LAST_ACCESS (0x00000020)
value FILE_NOTIFY_CHANGE_LAST_WRITE (0x00000010)
value FILE_NOTIFY_CHANGE_SECURITY (0x00000100)
value FILE_NOTIFY_CHANGE_SIZE (0x00000008)
value FILE_PERSISTENT_ACLS (0x00000008)
value FILE_PREFETCH_TYPE_FOR_CREATE (0x1)
value FILE_PREFETCH_TYPE_FOR_CREATE_EX (0x3)
value FILE_PREFETCH_TYPE_FOR_DIRENUM (0x2)
value FILE_PREFETCH_TYPE_FOR_DIRENUM_EX (0x4)
value FILE_PREFETCH_TYPE_MAX (0x4)
value FILE_PROVIDER_COMPRESSION_LZX ((0x00000001))
value FILE_PROVIDER_COMPRESSION_MAXIMUM ((0x00000004))
value FILE_PROVIDER_CURRENT_VERSION ((0x00000001))
value FILE_PROVIDER_FLAG_COMPRESS_ON_WRITE ((0x00000001))
value FILE_PROVIDER_SINGLE_FILE ((0x00000001))
value FILE_READ_ACCESS (( 0x0001 ))
value FILE_READ_ATTRIBUTES (( 0x0080 ))
value FILE_READ_DATA (( 0x0001 ))
value FILE_READ_EA (( 0x0008 ))
value FILE_READ_ONLY (8)
value FILE_READ_ONLY_VOLUME (0x00080000)
value FILE_REGION_USAGE_HUGE_PAGE_ALIGNMENT (0x00000010)
value FILE_REGION_USAGE_LARGE_PAGE_ALIGNMENT (0x00000008)
value FILE_REGION_USAGE_OTHER_PAGE_ALIGNMENT (0x00000004)
value FILE_REGION_USAGE_QUERY_ALIGNMENT ((FILE_REGION_USAGE_LARGE_PAGE_ALIGNMENT | FILE_REGION_USAGE_HUGE_PAGE_ALIGNMENT))
value FILE_REGION_USAGE_VALID_CACHED_DATA (0x00000001)
value FILE_REGION_USAGE_VALID_NONCACHED_DATA (0x00000002)
value FILE_RENAME_FLAG_POSIX_SEMANTICS (0x00000002)
value FILE_RENAME_FLAG_REPLACE_IF_EXISTS (0x00000001)
value FILE_RENAME_FLAG_SUPPRESS_PIN_STATE_INHERITANCE (0x00000004)
value FILE_RETURNS_CLEANUP_RESULT_INFO (0x00000200)
value FILE_ROOT_DIR (3)
value FILE_SEQUENTIAL_WRITE_ONCE (0x00100000)
value FILE_SET_ENCRYPTION (0x00000001)
value FILE_SHARE_DELETE (0x00000004)
value FILE_SHARE_READ (0x00000001)
value FILE_SHARE_WRITE (0x00000002)
value FILE_SKIP_COMPLETION_PORT_ON_SUCCESS (0x1)
value FILE_SKIP_SET_EVENT_ON_HANDLE (0x2)
value FILE_SPECIAL_ACCESS ((FILE_ANY_ACCESS))
value FILE_STORAGE_TIER_DESCRIPTION_LENGTH ((512))
value FILE_STORAGE_TIER_FLAG_NO_SEEK_PENALTY ((0x00020000))
value FILE_STORAGE_TIER_FLAG_PARITY ((0x00800000))
value FILE_STORAGE_TIER_FLAG_READ_CACHE ((0x00400000))
value FILE_STORAGE_TIER_FLAG_SMR ((0x01000000))
value FILE_STORAGE_TIER_FLAG_WRITE_BACK_CACHE ((0x00200000))
value FILE_STORAGE_TIER_NAME_LENGTH ((256))
value FILE_SUPPORTS_BLOCK_REFCOUNTING (0x08000000)
value FILE_SUPPORTS_BYPASS_IO (0x00000800)
value FILE_SUPPORTS_CASE_SENSITIVE_DIRS (0x00002000)
value FILE_SUPPORTS_ENCRYPTION (0x00020000)
value FILE_SUPPORTS_EXTENDED_ATTRIBUTES (0x00800000)
value FILE_SUPPORTS_GHOSTING (0x40000000)
value FILE_SUPPORTS_HARD_LINKS (0x00400000)
value FILE_SUPPORTS_INTEGRITY_STREAMS (0x04000000)
value FILE_SUPPORTS_OBJECT_IDS (0x00010000)
value FILE_SUPPORTS_OPEN_BY_FILE_ID (0x01000000)
value FILE_SUPPORTS_POSIX_UNLINK_RENAME (0x00000400)
value FILE_SUPPORTS_REMOTE_STORAGE (0x00000100)
value FILE_SUPPORTS_REPARSE_POINTS (0x00000080)
value FILE_SUPPORTS_SPARSE_FILES (0x00000040)
value FILE_SUPPORTS_SPARSE_VDL (0x10000000)
value FILE_SUPPORTS_STREAM_SNAPSHOTS (0x00001000)
value FILE_SUPPORTS_TRANSACTIONS (0x00200000)
value FILE_SUPPORTS_USN_JOURNAL (0x02000000)
value FILE_SYSTEM_ATTR (2)
value FILE_SYSTEM_DIR (4)
value FILE_SYSTEM_NOT_SUPPORT (6)
value FILE_TRAVERSE (( 0x0020 ))
value FILE_TYPE_CHAR (0x0002)
value FILE_TYPE_DISK (0x0001)
value FILE_TYPE_NOTIFICATION_FLAG_USAGE_BEGIN (0x00000001)
value FILE_TYPE_NOTIFICATION_FLAG_USAGE_END (0x00000002)
value FILE_TYPE_PIPE (0x0003)
value FILE_TYPE_REMOTE (0x8000)
value FILE_TYPE_UNKNOWN (0x0000)
value FILE_UNICODE_ON_DISK (0x00000004)
value FILE_UNKNOWN (5)
value FILE_USER_DISALLOWED (7)
value FILE_VER_GET_LOCALISED (0x01)
value FILE_VER_GET_NEUTRAL (0x02)
value FILE_VER_GET_PREFETCHED (0x04)
value FILE_VOLUME_IS_COMPRESSED (0x00008000)
value FILE_VOLUME_QUOTAS (0x00000020)
value FILE_WRITE_ACCESS (( 0x0002 ))
value FILE_WRITE_ATTRIBUTES (( 0x0100 ))
value FILE_WRITE_DATA (( 0x0002 ))
value FILE_WRITE_EA (( 0x0010 ))
value FILE_ZERO_DATA_INFORMATION_FLAG_PRESERVE_CACHED_DATA ((0x00000001))
value FILL_NV_MEMORY_FLAG_FLUSH ((0x00000001))
value FILL_NV_MEMORY_FLAG_NON_TEMPORAL ((0x00000002))
value FILL_NV_MEMORY_FLAG_NO_DRAIN ((0x00000100))
value FILL_NV_MEMORY_FLAG_PERSIST ((FILL_NV_MEMORY_FLAG_FLUSH | FILL_NV_MEMORY_FLAG_NON_TEMPORAL))
value FINDDLGORD (1540)
value FINDMSGSTRING (FINDMSGSTRINGA)
value FIND_ACTCTX_SECTION_KEY_RETURN_ASSEMBLY_METADATA ((0x00000004))
value FIND_ACTCTX_SECTION_KEY_RETURN_FLAGS ((0x00000002))
value FIND_ACTCTX_SECTION_KEY_RETURN_HACTCTX ((0x00000001))
value FIND_ENDSWITH (0x00200000)
value FIND_FIRST_EX_CASE_SENSITIVE (0x00000001)
value FIND_FIRST_EX_LARGE_FETCH (0x00000002)
value FIND_FIRST_EX_ON_DISK_ENTRIES_ONLY (0x00000004)
value FIND_FROMEND (0x00800000)
value FIND_FROMSTART (0x00400000)
value FIND_RESOURCE_DIRECTORY_LANGUAGES ((0x0400))
value FIND_RESOURCE_DIRECTORY_NAMES ((0x0200))
value FIND_RESOURCE_DIRECTORY_TYPES ((0x0100))
value FIND_STARTSWITH (0x00100000)
value FIXED_PITCH (1)
value FKF_AVAILABLE (0x00000002)
value FKF_CLICKON (0x00000040)
value FKF_CONFIRMHOTKEY (0x00000008)
value FKF_FILTERKEYSON (0x00000001)
value FKF_HOTKEYACTIVE (0x00000004)
value FKF_HOTKEYSOUND (0x00000010)
value FKF_INDICATOR (0x00000020)
value FLAG_USN_TRACK_MODIFIED_RANGES_ENABLE (0x00000001)
value FLASHW_ALL ((FLASHW_CAPTION | FLASHW_TRAY))
value FLASHW_CAPTION (0x00000001)
value FLASHW_STOP (0)
value FLASHW_TIMER (0x00000004)
value FLASHW_TIMERNOFG (0x0000000C)
value FLASHW_TRAY (0x00000002)
value FLI_GLYPHS (0x00040000L)
value FLI_MASK (0x103B)
value FLOODFILLBORDER (0)
value FLOODFILLSURFACE (1)
value FLS_MAXIMUM_AVAILABLE (4080)
value FLS_OUT_OF_INDEXES (((DWORD)0xFFFFFFFF))
value FLUSHOUTPUT (6)
value FLUSH_FLAGS_FILE_DATA_ONLY (0x00000001)
value FLUSH_FLAGS_FILE_DATA_SYNC_ONLY (0x00000004)
value FLUSH_FLAGS_NO_SYNC (0x00000002)
value FLUSH_NV_MEMORY_DEFAULT_TOKEN ((ULONG_PTR)(-1))
value FLUSH_NV_MEMORY_IN_FLAG_NO_DRAIN ((0x00000001))
value FMFD_DEFAULT (0x00000000)
value FMFD_ENABLEMIMESNIFFING (0x00000002)
value FMFD_IGNOREMIMETEXTPLAIN (0x00000004)
value FMFD_RESPECTTEXTPLAIN (0x00000010)
value FMFD_RETURNUPDATEDIMGMIMES (0x00000020)
value FMFD_SERVERMIME (0x00000008)
value FMFD_URLASFILENAME (0x00000001)
value FMTID_NULL (GUID_NULL)
value FNERR_BUFFERTOOSMALL (0x3003)
value FNERR_FILENAMECODES (0x3000)
value FNERR_INVALIDFILENAME (0x3002)
value FNERR_SUBCLASSFAILURE (0x3001)
value FNOINVERT (0x02)
value FOCUS_EVENT (0x0010)
value FOF_ALLOWUNDO (0x0040)
value FOF_CONFIRMMOUSE (0x0002)
value FOF_FILESONLY (0x0080)
value FOF_MULTIDESTFILES (0x0001)
value FOF_NOCONFIRMATION (0x0010)
value FOF_NOCONFIRMMKDIR (0x0200)
value FOF_NOCOPYSECURITYATTRIBS (0x0800)
value FOF_NOERRORUI (0x0400)
value FOF_NORECURSEREPARSE (0x8000)
value FOF_NORECURSION (0x1000)
value FOF_NO_CONNECTED_ELEMENTS (0x2000)
value FOF_NO_UI ((FOF_SILENT | FOF_NOCONFIRMATION | FOF_NOERRORUI | FOF_NOCONFIRMMKDIR))
value FOF_RENAMEONCOLLISION (0x0008)
value FOF_SILENT (0x0004)
value FOF_SIMPLEPROGRESS (0x0100)
value FOF_WANTMAPPINGHANDLE (0x0020)
value FOF_WANTNUKEWARNING (0x4000)
value FONTDLGORD (1542)
value FONTMAPPER_MAX (10)
value FOPEN_MAX (20)
value FOREGROUND_BLUE (0x0001)
value FOREGROUND_GREEN (0x0002)
value FOREGROUND_INTENSITY (0x0008)
value FOREGROUND_RED (0x0004)
value FOREST_USER_RID_MAX ((0x000001F3L))
value FORMAT_MESSAGE_ALLOCATE_BUFFER (0x00000100)
value FORMAT_MESSAGE_ARGUMENT_ARRAY (0x00002000)
value FORMAT_MESSAGE_FROM_HMODULE (0x00000800)
value FORMAT_MESSAGE_FROM_STRING (0x00000400)
value FORMAT_MESSAGE_FROM_SYSTEM (0x00001000)
value FORMAT_MESSAGE_IGNORE_INSERTS (0x00000200)
value FORMAT_MESSAGE_MAX_WIDTH_MASK (0x000000FF)
value FORM_BUILTIN (0x00000001)
value FORM_PRINTER (0x00000002)
value FORM_USER (0x00000000)
value FO_COPY (0x0002)
value FO_DELETE (0x0003)
value FO_MOVE (0x0001)
value FO_RENAME (0x0004)
value FRAME_FPO (0)
value FRAME_NONFPO (3)
value FRAME_TRAP (1)
value FRAME_TSS (2)
value FRERR_BUFFERLENGTHZERO (0x4001)
value FRERR_FINDREPLACECODES (0x4000)
value FRM_FIRST ((WM_USER + 100))
value FRM_LAST ((WM_USER + 200))
value FRM_SETOPERATIONRESULT ((FRM_FIRST + 0x0000))
value FRM_SETOPERATIONRESULTTEXT ((FRM_FIRST + 0x0001))
value FROM_PROTOCOL_INFO ((-1))
value FRS_ERR_AUTHENTICATION (8008)
value FRS_ERR_CHILD_TO_PARENT_COMM (8011)
value FRS_ERR_INSUFFICIENT_PRIV (8007)
value FRS_ERR_INTERNAL (8005)
value FRS_ERR_INTERNAL_API (8004)
value FRS_ERR_INVALID_API_SEQUENCE (8001)
value FRS_ERR_INVALID_SERVICE_PARAMETER (8017)
value FRS_ERR_PARENT_AUTHENTICATION (8010)
value FRS_ERR_PARENT_INSUFFICIENT_PRIV (8009)
value FRS_ERR_PARENT_TO_CHILD_COMM (8012)
value FRS_ERR_SERVICE_COMM (8006)
value FRS_ERR_STARTING_SERVICE (8002)
value FRS_ERR_STOPPING_SERVICE (8003)
value FRS_ERR_SYSVOL_DEMOTE (8016)
value FRS_ERR_SYSVOL_IS_BUSY (8015)
value FRS_ERR_SYSVOL_POPULATE (8013)
value FRS_ERR_SYSVOL_POPULATE_TIMEOUT (8014)
value FR_DIALOGTERM (0x00000040)
value FR_DOWN (0x00000001)
value FR_ENABLEHOOK (0x00000100)
value FR_ENABLETEMPLATE (0x00000200)
value FR_ENABLETEMPLATEHANDLE (0x00002000)
value FR_FINDNEXT (0x00000008)
value FR_HIDEMATCHCASE (0x00008000)
value FR_HIDEUPDOWN (0x00004000)
value FR_HIDEWHOLEWORD (0x00010000)
value FR_MATCHALEFHAMZA (0x80000000)
value FR_MATCHCASE (0x00000004)
value FR_MATCHDIAC (0x20000000)
value FR_MATCHKASHIDA (0x40000000)
value FR_NOMATCHCASE (0x00000800)
value FR_NOT_ENUM (0x20)
value FR_NOUPDOWN (0x00000400)
value FR_NOWHOLEWORD (0x00001000)
value FR_NOWRAPAROUND (0x00080000)
value FR_PRIVATE (0x10)
value FR_RAW (0x00020000)
value FR_REPLACE (0x00000010)
value FR_REPLACEALL (0x00000020)
value FR_SHOWHELP (0x00000080)
value FR_SHOWWRAPAROUND (0x00040000)
value FR_WHOLEWORD (0x00000002)
value FR_WRAPAROUND (0x00100000)
value FSCTL_INTEGRITY_FLAG_CHECKSUM_ENFORCEMENT_OFF ((1))
value FSCTL_MARK_AS_SYSTEM_HIVE (FSCTL_SET_BOOTLOADER_ACCESSED)
value FSHIFT (0x04)
value FS_ARABIC (0x00000040L)
value FS_BALTIC (0x00000080L)
value FS_CASE_IS_PRESERVED (FILE_CASE_PRESERVED_NAMES)
value FS_CASE_SENSITIVE (FILE_CASE_SENSITIVE_SEARCH)
value FS_CHINESESIMP (0x00040000L)
value FS_CHINESETRAD (0x00100000L)
value FS_CYRILLIC (0x00000004L)
value FS_FILE_COMPRESSION (FILE_FILE_COMPRESSION)
value FS_FILE_ENCRYPTION (FILE_SUPPORTS_ENCRYPTION)
value FS_GREEK (0x00000008L)
value FS_HEBREW (0x00000020L)
value FS_JISJAPAN (0x00020000L)
value FS_JOHAB (0x00200000L)
value FS_PERSISTENT_ACLS (FILE_PERSISTENT_ACLS)
value FS_SYMBOL (0x80000000L)
value FS_THAI (0x00010000L)
value FS_TURKISH (0x00000010L)
value FS_UNICODE_STORED_ON_DISK (FILE_UNICODE_ON_DISK)
value FS_VIETNAMESE (0x00000100L)
value FS_VOL_IS_COMPRESSED (FILE_VOLUME_IS_COMPRESSED)
value FS_WANSUNG (0x00080000L)
value FVE_E_AAD_ENDPOINT_BUSY (_HRESULT_TYPEDEF_(0x803100E1L))
value FVE_E_AAD_SERVER_FAIL_BACKOFF (_HRESULT_TYPEDEF_(0x803100EAL))
value FVE_E_AAD_SERVER_FAIL_RETRY_AFTER (_HRESULT_TYPEDEF_(0x803100E9L))
value FVE_E_ACTION_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310009L))
value FVE_E_ADBACKUP_NOT_ENABLED (_HRESULT_TYPEDEF_(0x803100D5L))
value FVE_E_AD_ATTR_NOT_SET (_HRESULT_TYPEDEF_(0x8031000EL))
value FVE_E_AD_BACKUP_REQUIRED_POLICY_NOT_SET_FIXED_DRIVE (_HRESULT_TYPEDEF_(0x803100DBL))
value FVE_E_AD_BACKUP_REQUIRED_POLICY_NOT_SET_OS_DRIVE (_HRESULT_TYPEDEF_(0x803100DAL))
value FVE_E_AD_BACKUP_REQUIRED_POLICY_NOT_SET_REMOVABLE_DRIVE (_HRESULT_TYPEDEF_(0x803100DCL))
value FVE_E_AD_GUID_NOT_FOUND (_HRESULT_TYPEDEF_(0x8031000FL))
value FVE_E_AD_INSUFFICIENT_BUFFER (_HRESULT_TYPEDEF_(0x8031001AL))
value FVE_E_AD_INVALID_DATASIZE (_HRESULT_TYPEDEF_(0x8031000CL))
value FVE_E_AD_INVALID_DATATYPE (_HRESULT_TYPEDEF_(0x8031000BL))
value FVE_E_AD_NO_VALUES (_HRESULT_TYPEDEF_(0x8031000DL))
value FVE_E_AD_SCHEMA_NOT_INSTALLED (_HRESULT_TYPEDEF_(0x8031000AL))
value FVE_E_AUTH_INVALID_APPLICATION (_HRESULT_TYPEDEF_(0x80310044L))
value FVE_E_AUTH_INVALID_CONFIG (_HRESULT_TYPEDEF_(0x80310045L))
value FVE_E_AUTOUNLOCK_ENABLED (_HRESULT_TYPEDEF_(0x80310029L))
value FVE_E_BAD_DATA (_HRESULT_TYPEDEF_(0x80310016L))
value FVE_E_BAD_INFORMATION (_HRESULT_TYPEDEF_(0x80310010L))
value FVE_E_BAD_PARTITION_SIZE (_HRESULT_TYPEDEF_(0x80310014L))
value FVE_E_BCD_APPLICATIONS_PATH_INCORRECT (_HRESULT_TYPEDEF_(0x80310052L))
value FVE_E_BOOTABLE_CDDVD (_HRESULT_TYPEDEF_(0x80310030L))
value FVE_E_BUFFER_TOO_LARGE (_HRESULT_TYPEDEF_(0x803100CFL))
value FVE_E_CANNOT_ENCRYPT_NO_KEY (_HRESULT_TYPEDEF_(0x8031002EL))
value FVE_E_CANNOT_SET_FVEK_ENCRYPTED (_HRESULT_TYPEDEF_(0x8031002DL))
value FVE_E_CANT_LOCK_AUTOUNLOCK_ENABLED_VOLUME (_HRESULT_TYPEDEF_(0x80310097L))
value FVE_E_CLUSTERING_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8031001EL))
value FVE_E_CONV_READ (_HRESULT_TYPEDEF_(0x8031001BL))
value FVE_E_CONV_RECOVERY_FAILED (_HRESULT_TYPEDEF_(0x80310088L))
value FVE_E_CONV_WRITE (_HRESULT_TYPEDEF_(0x8031001CL))
value FVE_E_DATASET_FULL (_HRESULT_TYPEDEF_(0x803100EBL))
value FVE_E_DEBUGGER_ENABLED (_HRESULT_TYPEDEF_(0x8031004FL))
value FVE_E_DEVICELOCKOUT_COUNTER_MISMATCH (_HRESULT_TYPEDEF_(0x803100CEL))
value FVE_E_DEVICE_LOCKOUT_COUNTER_UNAVAILABLE (_HRESULT_TYPEDEF_(0x803100CDL))
value FVE_E_DEVICE_NOT_JOINED (_HRESULT_TYPEDEF_(0x803100E0L))
value FVE_E_DE_DEVICE_LOCKEDOUT (_HRESULT_TYPEDEF_(0x803100CAL))
value FVE_E_DE_FIXED_DATA_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803100C5L))
value FVE_E_DE_HARDWARE_NOT_COMPLIANT (_HRESULT_TYPEDEF_(0x803100C6L))
value FVE_E_DE_OS_VOLUME_NOT_PROTECTED (_HRESULT_TYPEDEF_(0x803100C9L))
value FVE_E_DE_PREVENTED_FOR_OS (_HRESULT_TYPEDEF_(0x803100D1L))
value FVE_E_DE_PROTECTION_NOT_YET_ENABLED (_HRESULT_TYPEDEF_(0x803100CBL))
value FVE_E_DE_PROTECTION_SUSPENDED (_HRESULT_TYPEDEF_(0x803100C8L))
value FVE_E_DE_VOLUME_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803100D3L))
value FVE_E_DE_VOLUME_OPTED_OUT (_HRESULT_TYPEDEF_(0x803100D2L))
value FVE_E_DE_WINRE_NOT_CONFIGURED (_HRESULT_TYPEDEF_(0x803100C7L))
value FVE_E_DRY_RUN_FAILED (_HRESULT_TYPEDEF_(0x8031004DL))
value FVE_E_DV_NOT_ALLOWED_BY_GP (_HRESULT_TYPEDEF_(0x80310071L))
value FVE_E_DV_NOT_SUPPORTED_ON_FS (_HRESULT_TYPEDEF_(0x80310070L))
value FVE_E_EDRIVE_BAND_ENUMERATION_FAILED (_HRESULT_TYPEDEF_(0x803100E3L))
value FVE_E_EDRIVE_BAND_IN_USE (_HRESULT_TYPEDEF_(0x803100B0L))
value FVE_E_EDRIVE_DISALLOWED_BY_GP (_HRESULT_TYPEDEF_(0x803100B1L))
value FVE_E_EDRIVE_DRY_RUN_FAILED (_HRESULT_TYPEDEF_(0x803100BCL))
value FVE_E_EDRIVE_DV_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803100B4L))
value FVE_E_EDRIVE_INCOMPATIBLE_FIRMWARE (_HRESULT_TYPEDEF_(0x803100BFL))
value FVE_E_EDRIVE_INCOMPATIBLE_VOLUME (_HRESULT_TYPEDEF_(0x803100B2L))
value FVE_E_EDRIVE_NO_FAILOVER_TO_SW (_HRESULT_TYPEDEF_(0x803100AFL))
value FVE_E_EFI_ONLY (_HRESULT_TYPEDEF_(0x8031009CL))
value FVE_E_ENH_PIN_INVALID (_HRESULT_TYPEDEF_(0x80310099L))
value FVE_E_EOW_NOT_SUPPORTED_IN_VERSION (_HRESULT_TYPEDEF_(0x803100D4L))
value FVE_E_EXECUTE_REQUEST_SENT_TOO_SOON (_HRESULT_TYPEDEF_(0x803100DEL))
value FVE_E_FAILED_AUTHENTICATION (_HRESULT_TYPEDEF_(0x80310027L))
value FVE_E_FAILED_SECTOR_SIZE (_HRESULT_TYPEDEF_(0x80310026L))
value FVE_E_FAILED_WRONG_FS (_HRESULT_TYPEDEF_(0x80310013L))
value FVE_E_FIPS_DISABLE_PROTECTION_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310046L))
value FVE_E_FIPS_HASH_KDF_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310098L))
value FVE_E_FIPS_PREVENTS_EXTERNAL_KEY_EXPORT (_HRESULT_TYPEDEF_(0x80310038L))
value FVE_E_FIPS_PREVENTS_PASSPHRASE (_HRESULT_TYPEDEF_(0x8031006CL))
value FVE_E_FIPS_PREVENTS_RECOVERY_PASSWORD (_HRESULT_TYPEDEF_(0x80310037L))
value FVE_E_FIPS_RNG_CHECK_FAILED (_HRESULT_TYPEDEF_(0x80310036L))
value FVE_E_FIRMWARE_TYPE_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80310048L))
value FVE_E_FOREIGN_VOLUME (_HRESULT_TYPEDEF_(0x80310023L))
value FVE_E_FS_MOUNTED (_HRESULT_TYPEDEF_(0x8031004BL))
value FVE_E_FS_NOT_EXTENDED (_HRESULT_TYPEDEF_(0x80310047L))
value FVE_E_FULL_ENCRYPTION_NOT_ALLOWED_ON_TP_STORAGE (_HRESULT_TYPEDEF_(0x803100A5L))
value FVE_E_HIDDEN_VOLUME (_HRESULT_TYPEDEF_(0x80310056L))
value FVE_E_INVALID_BITLOCKER_OID (_HRESULT_TYPEDEF_(0x8031006EL))
value FVE_E_INVALID_DATUM_TYPE (_HRESULT_TYPEDEF_(0x8031009BL))
value FVE_E_INVALID_KEY_FORMAT (_HRESULT_TYPEDEF_(0x80310034L))
value FVE_E_INVALID_NBP_CERT (_HRESULT_TYPEDEF_(0x803100E2L))
value FVE_E_INVALID_NKP_CERT (_HRESULT_TYPEDEF_(0x8031009FL))
value FVE_E_INVALID_PASSWORD_FORMAT (_HRESULT_TYPEDEF_(0x80310035L))
value FVE_E_INVALID_PIN_CHARS (_HRESULT_TYPEDEF_(0x8031009AL))
value FVE_E_INVALID_PIN_CHARS_DETAILED (_HRESULT_TYPEDEF_(0x803100CCL))
value FVE_E_INVALID_PROTECTOR_TYPE (_HRESULT_TYPEDEF_(0x8031003AL))
value FVE_E_INVALID_STARTUP_OPTIONS (_HRESULT_TYPEDEF_(0x8031005BL))
value FVE_E_KEYFILE_INVALID (_HRESULT_TYPEDEF_(0x8031003DL))
value FVE_E_KEYFILE_NOT_FOUND (_HRESULT_TYPEDEF_(0x8031003CL))
value FVE_E_KEYFILE_NO_VMK (_HRESULT_TYPEDEF_(0x8031003EL))
value FVE_E_KEY_LENGTH_NOT_SUPPORTED_BY_EDRIVE (_HRESULT_TYPEDEF_(0x803100A7L))
value FVE_E_KEY_PROTECTOR_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80310069L))
value FVE_E_KEY_REQUIRED (_HRESULT_TYPEDEF_(0x8031001DL))
value FVE_E_KEY_ROTATION_NOT_ENABLED (_HRESULT_TYPEDEF_(0x803100DFL))
value FVE_E_KEY_ROTATION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803100DDL))
value FVE_E_LIVEID_ACCOUNT_BLOCKED (_HRESULT_TYPEDEF_(0x803100C3L))
value FVE_E_LIVEID_ACCOUNT_SUSPENDED (_HRESULT_TYPEDEF_(0x803100C2L))
value FVE_E_LOCKED_VOLUME (_HRESULT_TYPEDEF_(0x80310000L))
value FVE_E_METADATA_FULL (_HRESULT_TYPEDEF_(0x803100ECL))
value FVE_E_MOR_FAILED (_HRESULT_TYPEDEF_(0x80310055L))
value FVE_E_MULTIPLE_NKP_CERTS (_HRESULT_TYPEDEF_(0x8031009DL))
value FVE_E_NON_BITLOCKER_KU (_HRESULT_TYPEDEF_(0x80310093L))
value FVE_E_NON_BITLOCKER_OID (_HRESULT_TYPEDEF_(0x80310085L))
value FVE_E_NOT_ACTIVATED (_HRESULT_TYPEDEF_(0x80310008L))
value FVE_E_NOT_ALLOWED_IN_SAFE_MODE (_HRESULT_TYPEDEF_(0x80310040L))
value FVE_E_NOT_ALLOWED_IN_VERSION (_HRESULT_TYPEDEF_(0x80310053L))
value FVE_E_NOT_ALLOWED_ON_CLUSTER (_HRESULT_TYPEDEF_(0x803100AEL))
value FVE_E_NOT_ALLOWED_ON_CSV_STACK (_HRESULT_TYPEDEF_(0x803100ADL))
value FVE_E_NOT_ALLOWED_TO_UPGRADE_WHILE_CONVERTING (_HRESULT_TYPEDEF_(0x803100B3L))
value FVE_E_NOT_DATA_VOLUME (_HRESULT_TYPEDEF_(0x80310019L))
value FVE_E_NOT_DECRYPTED (_HRESULT_TYPEDEF_(0x80310039L))
value FVE_E_NOT_DE_VOLUME (_HRESULT_TYPEDEF_(0x803100D7L))
value FVE_E_NOT_ENCRYPTED (_HRESULT_TYPEDEF_(0x80310001L))
value FVE_E_NOT_ON_STACK (_HRESULT_TYPEDEF_(0x8031004AL))
value FVE_E_NOT_OS_VOLUME (_HRESULT_TYPEDEF_(0x80310028L))
value FVE_E_NOT_PROVISIONED_ON_ALL_VOLUMES (_HRESULT_TYPEDEF_(0x803100C4L))
value FVE_E_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80310015L))
value FVE_E_NO_AUTOUNLOCK_MASTER_KEY (_HRESULT_TYPEDEF_(0x80310054L))
value FVE_E_NO_BOOTMGR_METRIC (_HRESULT_TYPEDEF_(0x80310005L))
value FVE_E_NO_BOOTSECTOR_METRIC (_HRESULT_TYPEDEF_(0x80310004L))
value FVE_E_NO_EXISTING_PASSPHRASE (_HRESULT_TYPEDEF_(0x803100A8L))
value FVE_E_NO_EXISTING_PIN (_HRESULT_TYPEDEF_(0x803100A0L))
value FVE_E_NO_FEATURE_LICENSE (_HRESULT_TYPEDEF_(0x8031005AL))
value FVE_E_NO_LICENSE (_HRESULT_TYPEDEF_(0x80310049L))
value FVE_E_NO_MBR_METRIC (_HRESULT_TYPEDEF_(0x80310003L))
value FVE_E_NO_PASSPHRASE_WITH_TPM (_HRESULT_TYPEDEF_(0x803100ABL))
value FVE_E_NO_PREBOOT_KEYBOARD_DETECTED (_HRESULT_TYPEDEF_(0x803100B5L))
value FVE_E_NO_PREBOOT_KEYBOARD_OR_WINRE_DETECTED (_HRESULT_TYPEDEF_(0x803100B6L))
value FVE_E_NO_PROTECTORS_TO_TEST (_HRESULT_TYPEDEF_(0x8031003BL))
value FVE_E_NO_SUCH_CAPABILITY_ON_TARGET (_HRESULT_TYPEDEF_(0x803100D0L))
value FVE_E_NO_TPM_BIOS (_HRESULT_TYPEDEF_(0x80310002L))
value FVE_E_NO_TPM_WITH_PASSPHRASE (_HRESULT_TYPEDEF_(0x803100ACL))
value FVE_E_OPERATION_NOT_SUPPORTED_ON_VISTA_VOLUME (_HRESULT_TYPEDEF_(0x80310096L))
value FVE_E_OSV_KSR_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x803100D9L))
value FVE_E_OS_NOT_PROTECTED (_HRESULT_TYPEDEF_(0x80310020L))
value FVE_E_OS_VOLUME_PASSPHRASE_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x8031006DL))
value FVE_E_OVERLAPPED_UPDATE (_HRESULT_TYPEDEF_(0x80310024L))
value FVE_E_PASSPHRASE_PROTECTOR_CHANGE_BY_STD_USER_DISALLOWED (_HRESULT_TYPEDEF_(0x803100C1L))
value FVE_E_PASSPHRASE_TOO_LONG (_HRESULT_TYPEDEF_(0x803100AAL))
value FVE_E_PIN_INVALID (_HRESULT_TYPEDEF_(0x80310043L))
value FVE_E_PIN_PROTECTOR_CHANGE_BY_STD_USER_DISALLOWED (_HRESULT_TYPEDEF_(0x803100A2L))
value FVE_E_POLICY_CONFLICT_FDV_RK_OFF_AUK_ON (_HRESULT_TYPEDEF_(0x80310083L))
value FVE_E_POLICY_CONFLICT_FDV_RP_OFF_ADB_ON (_HRESULT_TYPEDEF_(0x80310091L))
value FVE_E_POLICY_CONFLICT_OSV_RP_OFF_ADB_ON (_HRESULT_TYPEDEF_(0x80310090L))
value FVE_E_POLICY_CONFLICT_RDV_RK_OFF_AUK_ON (_HRESULT_TYPEDEF_(0x80310084L))
value FVE_E_POLICY_CONFLICT_RDV_RP_OFF_ADB_ON (_HRESULT_TYPEDEF_(0x80310092L))
value FVE_E_POLICY_CONFLICT_RO_AND_STARTUP_KEY_REQUIRED (_HRESULT_TYPEDEF_(0x80310087L))
value FVE_E_POLICY_INVALID_ENHANCED_BCD_SETTINGS (_HRESULT_TYPEDEF_(0x803100BEL))
value FVE_E_POLICY_INVALID_PASSPHRASE_LENGTH (_HRESULT_TYPEDEF_(0x80310080L))
value FVE_E_POLICY_INVALID_PIN_LENGTH (_HRESULT_TYPEDEF_(0x80310068L))
value FVE_E_POLICY_ON_RDV_EXCLUSION_LIST (_HRESULT_TYPEDEF_(0x803100E4L))
value FVE_E_POLICY_PASSPHRASE_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x8031006AL))
value FVE_E_POLICY_PASSPHRASE_REQUIRED (_HRESULT_TYPEDEF_(0x8031006BL))
value FVE_E_POLICY_PASSPHRASE_REQUIRES_ASCII (_HRESULT_TYPEDEF_(0x803100A4L))
value FVE_E_POLICY_PASSPHRASE_TOO_SIMPLE (_HRESULT_TYPEDEF_(0x80310081L))
value FVE_E_POLICY_PASSWORD_REQUIRED (_HRESULT_TYPEDEF_(0x8031002CL))
value FVE_E_POLICY_PROHIBITS_SELFSIGNED (_HRESULT_TYPEDEF_(0x80310086L))
value FVE_E_POLICY_RECOVERY_KEY_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x8031005EL))
value FVE_E_POLICY_RECOVERY_KEY_REQUIRED (_HRESULT_TYPEDEF_(0x8031005FL))
value FVE_E_POLICY_RECOVERY_PASSWORD_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x8031005CL))
value FVE_E_POLICY_RECOVERY_PASSWORD_REQUIRED (_HRESULT_TYPEDEF_(0x8031005DL))
value FVE_E_POLICY_REQUIRES_RECOVERY_PASSWORD_ON_TOUCH_DEVICE (_HRESULT_TYPEDEF_(0x803100B8L))
value FVE_E_POLICY_REQUIRES_STARTUP_PIN_ON_TOUCH_DEVICE (_HRESULT_TYPEDEF_(0x803100B7L))
value FVE_E_POLICY_STARTUP_KEY_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310062L))
value FVE_E_POLICY_STARTUP_KEY_REQUIRED (_HRESULT_TYPEDEF_(0x80310063L))
value FVE_E_POLICY_STARTUP_PIN_KEY_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310064L))
value FVE_E_POLICY_STARTUP_PIN_KEY_REQUIRED (_HRESULT_TYPEDEF_(0x80310065L))
value FVE_E_POLICY_STARTUP_PIN_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310060L))
value FVE_E_POLICY_STARTUP_PIN_REQUIRED (_HRESULT_TYPEDEF_(0x80310061L))
value FVE_E_POLICY_STARTUP_TPM_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310066L))
value FVE_E_POLICY_STARTUP_TPM_REQUIRED (_HRESULT_TYPEDEF_(0x80310067L))
value FVE_E_POLICY_USER_CERTIFICATE_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310072L))
value FVE_E_POLICY_USER_CERTIFICATE_REQUIRED (_HRESULT_TYPEDEF_(0x80310073L))
value FVE_E_POLICY_USER_CERT_MUST_BE_HW (_HRESULT_TYPEDEF_(0x80310074L))
value FVE_E_POLICY_USER_CONFIGURE_FDV_AUTOUNLOCK_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310075L))
value FVE_E_POLICY_USER_CONFIGURE_RDV_AUTOUNLOCK_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310076L))
value FVE_E_POLICY_USER_CONFIGURE_RDV_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310077L))
value FVE_E_POLICY_USER_DISABLE_RDV_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310079L))
value FVE_E_POLICY_USER_ENABLE_RDV_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310078L))
value FVE_E_PREDICTED_TPM_PROTECTOR_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803100E5L))
value FVE_E_PRIVATEKEY_AUTH_FAILED (_HRESULT_TYPEDEF_(0x80310094L))
value FVE_E_PROTECTION_CANNOT_BE_DISABLED (_HRESULT_TYPEDEF_(0x803100D8L))
value FVE_E_PROTECTION_DISABLED (_HRESULT_TYPEDEF_(0x80310021L))
value FVE_E_PROTECTOR_CHANGE_MAX_PASSPHRASE_CHANGE_ATTEMPTS_REACHED (_HRESULT_TYPEDEF_(0x803100C0L))
value FVE_E_PROTECTOR_CHANGE_MAX_PIN_CHANGE_ATTEMPTS_REACHED (_HRESULT_TYPEDEF_(0x803100A3L))
value FVE_E_PROTECTOR_CHANGE_PASSPHRASE_MISMATCH (_HRESULT_TYPEDEF_(0x803100A9L))
value FVE_E_PROTECTOR_CHANGE_PIN_MISMATCH (_HRESULT_TYPEDEF_(0x803100A1L))
value FVE_E_PROTECTOR_EXISTS (_HRESULT_TYPEDEF_(0x80310031L))
value FVE_E_PROTECTOR_NOT_FOUND (_HRESULT_TYPEDEF_(0x80310033L))
value FVE_E_PUBKEY_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80310058L))
value FVE_E_RAW_ACCESS (_HRESULT_TYPEDEF_(0x80310050L))
value FVE_E_RAW_BLOCKED (_HRESULT_TYPEDEF_(0x80310051L))
value FVE_E_REBOOT_REQUIRED (_HRESULT_TYPEDEF_(0x8031004EL))
value FVE_E_RECOVERY_KEY_REQUIRED (_HRESULT_TYPEDEF_(0x80310022L))
value FVE_E_RECOVERY_PARTITION (_HRESULT_TYPEDEF_(0x80310082L))
value FVE_E_RELATIVE_PATH (_HRESULT_TYPEDEF_(0x80310032L))
value FVE_E_REMOVAL_OF_DRA_FAILED (_HRESULT_TYPEDEF_(0x80310095L))
value FVE_E_REMOVAL_OF_NKP_FAILED (_HRESULT_TYPEDEF_(0x8031009EL))
value FVE_E_SECUREBOOT_CONFIGURATION_INVALID (_HRESULT_TYPEDEF_(0x803100BBL))
value FVE_E_SECUREBOOT_DISABLED (_HRESULT_TYPEDEF_(0x803100BAL))
value FVE_E_SECURE_KEY_REQUIRED (_HRESULT_TYPEDEF_(0x80310007L))
value FVE_E_SETUP_TPM_CALLBACK_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803100E6L))
value FVE_E_SHADOW_COPY_PRESENT (_HRESULT_TYPEDEF_(0x803100BDL))
value FVE_E_SYSTEM_VOLUME (_HRESULT_TYPEDEF_(0x80310012L))
value FVE_E_TOKEN_NOT_IMPERSONATED (_HRESULT_TYPEDEF_(0x8031004CL))
value FVE_E_TOO_SMALL (_HRESULT_TYPEDEF_(0x80310011L))
value FVE_E_TPM_CONTEXT_SETUP_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803100E7L))
value FVE_E_TPM_DISABLED (_HRESULT_TYPEDEF_(0x8031003FL))
value FVE_E_TPM_INVALID_PCR (_HRESULT_TYPEDEF_(0x80310041L))
value FVE_E_TPM_NOT_OWNED (_HRESULT_TYPEDEF_(0x80310018L))
value FVE_E_TPM_NO_VMK (_HRESULT_TYPEDEF_(0x80310042L))
value FVE_E_TPM_SRK_AUTH_NOT_ZERO (_HRESULT_TYPEDEF_(0x80310025L))
value FVE_E_TRANSIENT_STATE (_HRESULT_TYPEDEF_(0x80310057L))
value FVE_E_UPDATE_INVALID_CONFIG (_HRESULT_TYPEDEF_(0x803100E8L))
value FVE_E_VIRTUALIZED_SPACE_TOO_BIG (_HRESULT_TYPEDEF_(0x80310089L))
value FVE_E_VOLUME_BOUND_ALREADY (_HRESULT_TYPEDEF_(0x8031001FL))
value FVE_E_VOLUME_EXTEND_PREVENTS_EOW_DECRYPT (_HRESULT_TYPEDEF_(0x803100D6L))
value FVE_E_VOLUME_HANDLE_OPEN (_HRESULT_TYPEDEF_(0x80310059L))
value FVE_E_VOLUME_NOT_BOUND (_HRESULT_TYPEDEF_(0x80310017L))
value FVE_E_VOLUME_TOO_SMALL (_HRESULT_TYPEDEF_(0x8031006FL))
value FVE_E_WIPE_CANCEL_NOT_APPLICABLE (_HRESULT_TYPEDEF_(0x803100B9L))
value FVE_E_WIPE_NOT_ALLOWED_ON_TP_STORAGE (_HRESULT_TYPEDEF_(0x803100A6L))
value FVE_E_WRONG_BOOTMGR (_HRESULT_TYPEDEF_(0x80310006L))
value FVE_E_WRONG_BOOTSECTOR (_HRESULT_TYPEDEF_(0x8031002AL))
value FVE_E_WRONG_SYSTEM_FS (_HRESULT_TYPEDEF_(0x8031002BL))
value FVIRTKEY (TRUE)
value FWP_E_ACTION_INCOMPATIBLE_WITH_LAYER (_HRESULT_TYPEDEF_(0x8032002CL))
value FWP_E_ACTION_INCOMPATIBLE_WITH_SUBLAYER (_HRESULT_TYPEDEF_(0x8032002DL))
value FWP_E_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x80320009L))
value FWP_E_BUILTIN_OBJECT (_HRESULT_TYPEDEF_(0x80320017L))
value FWP_E_CALLOUT_NOTIFICATION_FAILED (_HRESULT_TYPEDEF_(0x80320037L))
value FWP_E_CALLOUT_NOT_FOUND (_HRESULT_TYPEDEF_(0x80320001L))
value FWP_E_CONDITION_NOT_FOUND (_HRESULT_TYPEDEF_(0x80320002L))
value FWP_E_CONNECTIONS_DISABLED (_HRESULT_TYPEDEF_(0x80320041L))
value FWP_E_CONTEXT_INCOMPATIBLE_WITH_CALLOUT (_HRESULT_TYPEDEF_(0x8032002FL))
value FWP_E_CONTEXT_INCOMPATIBLE_WITH_LAYER (_HRESULT_TYPEDEF_(0x8032002EL))
value FWP_E_DROP_NOICMP (_HRESULT_TYPEDEF_(0x80320104L))
value FWP_E_DUPLICATE_AUTH_METHOD (_HRESULT_TYPEDEF_(0x8032003CL))
value FWP_E_DUPLICATE_CONDITION (_HRESULT_TYPEDEF_(0x8032002AL))
value FWP_E_DUPLICATE_KEYMOD (_HRESULT_TYPEDEF_(0x8032002BL))
value FWP_E_DYNAMIC_SESSION_IN_PROGRESS (_HRESULT_TYPEDEF_(0x8032000BL))
value FWP_E_EM_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80320032L))
value FWP_E_FILTER_NOT_FOUND (_HRESULT_TYPEDEF_(0x80320003L))
value FWP_E_IKEEXT_NOT_RUNNING (_HRESULT_TYPEDEF_(0x80320044L))
value FWP_E_INCOMPATIBLE_AUTH_METHOD (_HRESULT_TYPEDEF_(0x80320030L))
value FWP_E_INCOMPATIBLE_CIPHER_TRANSFORM (_HRESULT_TYPEDEF_(0x8032003AL))
value FWP_E_INCOMPATIBLE_DH_GROUP (_HRESULT_TYPEDEF_(0x80320031L))
value FWP_E_INCOMPATIBLE_LAYER (_HRESULT_TYPEDEF_(0x80320014L))
value FWP_E_INCOMPATIBLE_SA_STATE (_HRESULT_TYPEDEF_(0x8032001BL))
value FWP_E_INCOMPATIBLE_TXN (_HRESULT_TYPEDEF_(0x80320011L))
value FWP_E_INVALID_ACTION_TYPE (_HRESULT_TYPEDEF_(0x80320024L))
value FWP_E_INVALID_AUTH_TRANSFORM (_HRESULT_TYPEDEF_(0x80320038L))
value FWP_E_INVALID_CIPHER_TRANSFORM (_HRESULT_TYPEDEF_(0x80320039L))
value FWP_E_INVALID_DNS_NAME (_HRESULT_TYPEDEF_(0x80320042L))
value FWP_E_INVALID_ENUMERATOR (_HRESULT_TYPEDEF_(0x8032001DL))
value FWP_E_INVALID_FLAGS (_HRESULT_TYPEDEF_(0x8032001EL))
value FWP_E_INVALID_INTERVAL (_HRESULT_TYPEDEF_(0x80320021L))
value FWP_E_INVALID_NET_MASK (_HRESULT_TYPEDEF_(0x8032001FL))
value FWP_E_INVALID_PARAMETER (_HRESULT_TYPEDEF_(0x80320035L))
value FWP_E_INVALID_RANGE (_HRESULT_TYPEDEF_(0x80320020L))
value FWP_E_INVALID_TRANSFORM_COMBINATION (_HRESULT_TYPEDEF_(0x8032003BL))
value FWP_E_INVALID_TUNNEL_ENDPOINT (_HRESULT_TYPEDEF_(0x8032003DL))
value FWP_E_INVALID_WEIGHT (_HRESULT_TYPEDEF_(0x80320025L))
value FWP_E_IN_USE (_HRESULT_TYPEDEF_(0x8032000AL))
value FWP_E_KEY_DICTATION_INVALID_KEYING_MATERIAL (_HRESULT_TYPEDEF_(0x80320040L))
value FWP_E_KEY_DICTATOR_ALREADY_REGISTERED (_HRESULT_TYPEDEF_(0x8032003FL))
value FWP_E_KM_CLIENTS_ONLY (_HRESULT_TYPEDEF_(0x80320015L))
value FWP_E_LAYER_NOT_FOUND (_HRESULT_TYPEDEF_(0x80320004L))
value FWP_E_LIFETIME_MISMATCH (_HRESULT_TYPEDEF_(0x80320016L))
value FWP_E_MATCH_TYPE_MISMATCH (_HRESULT_TYPEDEF_(0x80320026L))
value FWP_E_NET_EVENTS_DISABLED (_HRESULT_TYPEDEF_(0x80320013L))
value FWP_E_NEVER_MATCH (_HRESULT_TYPEDEF_(0x80320033L))
value FWP_E_NOTIFICATION_DROPPED (_HRESULT_TYPEDEF_(0x80320019L))
value FWP_E_NOT_FOUND (_HRESULT_TYPEDEF_(0x80320008L))
value FWP_E_NO_TXN_IN_PROGRESS (_HRESULT_TYPEDEF_(0x8032000DL))
value FWP_E_NULL_DISPLAY_NAME (_HRESULT_TYPEDEF_(0x80320023L))
value FWP_E_NULL_POINTER (_HRESULT_TYPEDEF_(0x8032001CL))
value FWP_E_OUT_OF_BOUNDS (_HRESULT_TYPEDEF_(0x80320028L))
value FWP_E_PROVIDER_CONTEXT_MISMATCH (_HRESULT_TYPEDEF_(0x80320034L))
value FWP_E_PROVIDER_CONTEXT_NOT_FOUND (_HRESULT_TYPEDEF_(0x80320006L))
value FWP_E_PROVIDER_NOT_FOUND (_HRESULT_TYPEDEF_(0x80320005L))
value FWP_E_RESERVED (_HRESULT_TYPEDEF_(0x80320029L))
value FWP_E_SESSION_ABORTED (_HRESULT_TYPEDEF_(0x80320010L))
value FWP_E_STILL_ON (_HRESULT_TYPEDEF_(0x80320043L))
value FWP_E_SUBLAYER_NOT_FOUND (_HRESULT_TYPEDEF_(0x80320007L))
value FWP_E_TIMEOUT (_HRESULT_TYPEDEF_(0x80320012L))
value FWP_E_TOO_MANY_CALLOUTS (_HRESULT_TYPEDEF_(0x80320018L))
value FWP_E_TOO_MANY_SUBLAYERS (_HRESULT_TYPEDEF_(0x80320036L))
value FWP_E_TRAFFIC_MISMATCH (_HRESULT_TYPEDEF_(0x8032001AL))
value FWP_E_TXN_ABORTED (_HRESULT_TYPEDEF_(0x8032000FL))
value FWP_E_TXN_IN_PROGRESS (_HRESULT_TYPEDEF_(0x8032000EL))
value FWP_E_TYPE_MISMATCH (_HRESULT_TYPEDEF_(0x80320027L))
value FWP_E_WRONG_SESSION (_HRESULT_TYPEDEF_(0x8032000CL))
value FWP_E_ZERO_LENGTH_ARRAY (_HRESULT_TYPEDEF_(0x80320022L))
value FW_BLACK (FW_HEAVY)
value FW_BOLD (700)
value FW_DEMIBOLD (FW_SEMIBOLD)
value FW_DONTCARE (0)
value FW_EXTRABOLD (800)
value FW_EXTRALIGHT (200)
value FW_HEAVY (900)
value FW_ISSUEID_NO_ISSUE (0x00000000)
value FW_ISSUEID_UNKNOWN (0xFFFFFFFF)
value FW_LIGHT (300)
value FW_MEDIUM (500)
value FW_NORMAL (400)
value FW_REGULAR (FW_NORMAL)
value FW_SEMIBOLD (600)
value FW_THIN (100)
value FW_ULTRABOLD (FW_EXTRABOLD)
value FW_ULTRALIGHT (FW_EXTRALIGHT)
value GA_PARENT (1)
value GA_ROOT (2)
value GA_ROOTOWNER (3)
value GCF_INCLUDE_ANCESTORS (0x00000001)
value GCLP_HBRBACKGROUND ((-10))
value GCLP_HCURSOR ((-12))
value GCLP_HICON ((-14))
value GCLP_HICONSM ((-34))
value GCLP_HMODULE ((-16))
value GCLP_MENUNAME ((-8))
value GCLP_WNDPROC ((-24))
value GCL_CBCLSEXTRA ((-20))
value GCL_CBWNDEXTRA ((-18))
value GCL_CONVERSION (0x0001)
value GCL_REVERSECONVERSION (0x0002)
value GCL_REVERSE_LENGTH (0x0003)
value GCL_STYLE ((-26))
value GCN_E_DEFAULTNAMESPACE_EXISTS (_HRESULT_TYPEDEF_(0x803B0029L))
value GCN_E_MODULE_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0021L))
value GCN_E_NETADAPTER_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0026L))
value GCN_E_NETADAPTER_TIMEOUT (_HRESULT_TYPEDEF_(0x803B0025L))
value GCN_E_NETCOMPARTMENT_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0027L))
value GCN_E_NETINTERFACE_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0028L))
value GCN_E_NO_REQUEST_HANDLERS (_HRESULT_TYPEDEF_(0x803B0022L))
value GCN_E_REQUEST_UNSUPPORTED (_HRESULT_TYPEDEF_(0x803B0023L))
value GCN_E_RUNTIMEKEYS_FAILED (_HRESULT_TYPEDEF_(0x803B0024L))
value GCPCLASS_ARABIC (2)
value GCPCLASS_HEBREW (2)
value GCPCLASS_LATIN (1)
value GCPCLASS_LATINNUMBER (5)
value GCPCLASS_LATINNUMERICSEPARATOR (7)
value GCPCLASS_LATINNUMERICTERMINATOR (6)
value GCPCLASS_LOCALNUMBER (4)
value GCPCLASS_NEUTRAL (3)
value GCPCLASS_NUMERICSEPARATOR (8)
value GCPCLASS_POSTBOUNDLTR (0x20)
value GCPCLASS_POSTBOUNDRTL (0x10)
value GCPCLASS_PREBOUNDLTR (0x80)
value GCPCLASS_PREBOUNDRTL (0x40)
value GCPGLYPH_LINKAFTER (0x4000)
value GCPGLYPH_LINKBEFORE (0x8000)
value GCP_CLASSIN (0x00080000L)
value GCP_DBCS (0x0001)
value GCP_DIACRITIC (0x0100)
value GCP_DISPLAYZWG (0x00400000L)
value GCP_ERROR (0x8000)
value GCP_GLYPHSHAPE (0x0010)
value GCP_JUSTIFY (0x00010000L)
value GCP_JUSTIFYIN (0x00200000L)
value GCP_KASHIDA (0x0400)
value GCP_LIGATE (0x0020)
value GCP_MAXEXTENT (0x00100000L)
value GCP_NEUTRALOVERRIDE (0x02000000L)
value GCP_NUMERICOVERRIDE (0x01000000L)
value GCP_NUMERICSLATIN (0x04000000L)
value GCP_NUMERICSLOCAL (0x08000000L)
value GCP_REORDER (0x0002)
value GCP_SYMSWAPOFF (0x00800000L)
value GCP_USEKERNING (0x0008)
value GCS_COMPATTR (0x0010)
value GCS_COMPCLAUSE (0x0020)
value GCS_COMPREADATTR (0x0002)
value GCS_COMPREADCLAUSE (0x0004)
value GCS_COMPREADSTR (0x0001)
value GCS_COMPSTR (0x0008)
value GCS_CURSORPOS (0x0080)
value GCS_DELTASTART (0x0100)
value GCS_RESULTCLAUSE (0x1000)
value GCS_RESULTREADCLAUSE (0x0400)
value GCS_RESULTREADSTR (0x0200)
value GCS_RESULTSTR (0x0800)
value GCW_ATOM ((-32))
value GC_ALLGESTURES (0x00000001)
value GC_PAN (0x00000001)
value GC_PAN_WITH_GUTTER (0x00000008)
value GC_PAN_WITH_INERTIA (0x00000010)
value GC_PAN_WITH_SINGLE_FINGER_HORIZONTALLY (0x00000004)
value GC_PAN_WITH_SINGLE_FINGER_VERTICALLY (0x00000002)
value GC_PRESSANDTAP (0x00000001)
value GC_ROLLOVER (GC_PRESSANDTAP)
value GC_ROTATE (0x00000001)
value GC_TWOFINGERTAP (0x00000001)
value GC_ZOOM (0x00000001)
value GDICOMMENT_BEGINGROUP (0x00000002)
value GDICOMMENT_ENDGROUP (0x00000003)
value GDICOMMENT_IDENTIFIER (0x43494447)
value GDICOMMENT_MULTIFORMATS (0x40000004)
value GDICOMMENT_UNICODE_END (0x00000080)
value GDICOMMENT_UNICODE_STRING (0x00000040)
value GDICOMMENT_WINDOWS_METAFILE (0x80000001)
value GDIPLUS_TS_QUERYVER (4122)
value GDIPLUS_TS_RECORD (4123)
value GDI_ERROR ((0xFFFFFFFFL))
value GDI_MAX_OBJ_TYPE (GDI_OBJ_LAST)
value GDI_MIN_OBJ_TYPE (OBJ_PEN)
value GDI_OBJ_LAST (OBJ_COLORSPACE)
value GENERIC_ALL ((0x10000000L))
value GENERIC_EXECUTE ((0x20000000L))
value GENERIC_READ ((0x80000000L))
value GENERIC_WRITE ((0x40000000L))
value GEOID_NOT_AVAILABLE (-1)
value GEO_NAME_USER_DEFAULT (NULL)
value GESTURECONFIGMAXCOUNT (256)
value GESTUREVISUALIZATION_DOUBLETAP (0x0002)
value GESTUREVISUALIZATION_OFF (0x0000)
value GESTUREVISUALIZATION_ON (0x001F)
value GESTUREVISUALIZATION_PRESSANDHOLD (0x0008)
value GESTUREVISUALIZATION_PRESSANDTAP (0x0004)
value GESTUREVISUALIZATION_RIGHTTAP (0x0010)
value GESTUREVISUALIZATION_TAP (0x0001)
value GETCOLORTABLE (5)
value GETDEVICEUNITS (42)
value GETEXTENDEDTEXTMETRICS (256)
value GETEXTENTTABLE (257)
value GETFACENAME (513)
value GETPAIRKERNTABLE (258)
value GETPENWIDTH (16)
value GETPHYSPAGESIZE (12)
value GETPRINTINGOFFSET (13)
value GETSCALINGFACTOR (14)
value GETSETPAPERBINS (29)
value GETSETPAPERMETRICS (35)
value GETSETPRINTORIENT (30)
value GETSETSCREENPARAMS (3072)
value GETTECHNOLGY (20)
value GETTECHNOLOGY (20)
value GETTRACKKERNTABLE (259)
value GETVECTORBRUSHSIZE (27)
value GETVECTORPENSIZE (26)
value GET_FEATURE_FROM_PROCESS (0x00000002)
value GET_FEATURE_FROM_REGISTRY (0x00000004)
value GET_FEATURE_FROM_THREAD (0x00000001)
value GET_FEATURE_FROM_THREAD_INTERNET (0x00000040)
value GET_FEATURE_FROM_THREAD_INTRANET (0x00000010)
value GET_FEATURE_FROM_THREAD_LOCALMACHINE (0x00000008)
value GET_FEATURE_FROM_THREAD_RESTRICTED (0x00000080)
value GET_FEATURE_FROM_THREAD_TRUSTED (0x00000020)
value GET_MODULE_HANDLE_EX_FLAG_FROM_ADDRESS ((0x00000004))
value GET_MODULE_HANDLE_EX_FLAG_PIN ((0x00000001))
value GET_MODULE_HANDLE_EX_FLAG_UNCHANGED_REFCOUNT ((0x00000002))
value GET_MOUSEORKEY_LPARAM (GET_DEVICE_LPARAM)
value GET_PS_FEATURESETTING (4121)
value GET_TAPE_DRIVE_INFORMATION (1)
value GET_TAPE_MEDIA_INFORMATION (0)
value GET_VOLUME_BITMAP_FLAG_MASK_METADATA (0x00000001)
value GF_BEGIN (0x00000001)
value GF_END (0x00000004)
value GF_INERTIA (0x00000002)
value GGI_MARK_NONEXISTING_GLYPHS (0X0001)
value GGL_INDEX (0x00000002)
value GGL_LEVEL (0x00000001)
value GGL_PRIVATE (0x00000004)
value GGL_STRING (0x00000003)
value GGO_BEZIER (3)
value GGO_BITMAP (1)
value GGO_GLYPH_INDEX (0x0080)
value GGO_METRICS (0)
value GGO_NATIVE (2)
value GGO_UNHINTED (0x0100)
value GHND ((GMEM_MOVEABLE | GMEM_ZEROINIT))
value GIDC_ARRIVAL (1)
value GIDC_REMOVAL (2)
value GID_BEGIN (1)
value GID_END (2)
value GID_PAN (4)
value GID_PRESSANDTAP (7)
value GID_ROLLOVER (GID_PRESSANDTAP)
value GID_ROTATE (5)
value GID_TWOFINGERTAP (6)
value GID_ZOOM (3)
value GL_ID_CANNOTSAVE (0x00000011)
value GL_ID_CHOOSECANDIDATE (0x00000028)
value GL_ID_INPUTCODE (0x00000026)
value GL_ID_INPUTRADICAL (0x00000025)
value GL_ID_INPUTREADING (0x00000024)
value GL_ID_INPUTSYMBOL (0x00000027)
value GL_ID_NOCONVERT (0x00000020)
value GL_ID_NODICTIONARY (0x00000010)
value GL_ID_NOMODULE (0x00000001)
value GL_ID_PRIVATE_FIRST (0x00008000)
value GL_ID_PRIVATE_LAST (0x0000FFFF)
value GL_ID_READINGCONFLICT (0x00000023)
value GL_ID_REVERSECONVERSION (0x00000029)
value GL_ID_TOOMANYSTROKE (0x00000022)
value GL_ID_TYPINGERROR (0x00000021)
value GL_ID_UNKNOWN (0x00000000)
value GL_LEVEL_ERROR (0x00000002)
value GL_LEVEL_FATAL (0x00000001)
value GL_LEVEL_INFORMATION (0x00000004)
value GL_LEVEL_NOGUIDELINE (0x00000000)
value GL_LEVEL_WARNING (0x00000003)
value GMDI_GOINTOPOPUPS (0x0002L)
value GMDI_USEDISABLED (0x0001L)
value GMEM_DDESHARE (0x2000)
value GMEM_DISCARDABLE (0x0100)
value GMEM_DISCARDED (0x4000)
value GMEM_FIXED (0x0000)
value GMEM_INVALID_HANDLE (0x8000)
value GMEM_LOCKCOUNT (0x00FF)
value GMEM_LOWER (GMEM_NOT_BANKED)
value GMEM_MODIFY (0x0080)
value GMEM_MOVEABLE (0x0002)
value GMEM_NOCOMPACT (0x0010)
value GMEM_NODISCARD (0x0020)
value GMEM_NOTIFY (0x4000)
value GMEM_NOT_BANKED (0x1000)
value GMEM_SHARE (0x2000)
value GMEM_VALID_FLAGS (0x7F72)
value GMEM_ZEROINIT (0x0040)
value GMMP_USE_DISPLAY_POINTS (1)
value GMMP_USE_HIGH_RESOLUTION_POINTS (2)
value GM_ADVANCED (2)
value GM_COMPATIBLE (1)
value GM_LAST (2)
value GPTR ((GMEM_FIXED | GMEM_ZEROINIT))
value GPT_ATTRIBUTE_LEGACY_BIOS_BOOTABLE ((0x0000000000000004))
value GPT_ATTRIBUTE_NO_BLOCK_IO_PROTOCOL ((0x0000000000000002))
value GPT_ATTRIBUTE_PLATFORM_REQUIRED ((0x0000000000000001))
value GPT_BASIC_DATA_ATTRIBUTE_DAX ((0x0400000000000000))
value GPT_BASIC_DATA_ATTRIBUTE_HIDDEN ((0x4000000000000000))
value GPT_BASIC_DATA_ATTRIBUTE_NO_DRIVE_LETTER ((0x8000000000000000))
value GPT_BASIC_DATA_ATTRIBUTE_OFFLINE ((0x0800000000000000))
value GPT_BASIC_DATA_ATTRIBUTE_READ_ONLY ((0x1000000000000000))
value GPT_BASIC_DATA_ATTRIBUTE_SERVICE ((0x0200000000000000))
value GPT_BASIC_DATA_ATTRIBUTE_SHADOW_COPY ((0x2000000000000000))
value GPT_SPACES_ATTRIBUTE_NO_METADATA ((0x8000000000000000))
value GRADIENT_FILL_OP_FLAG (0x000000ff)
value GRADIENT_FILL_RECT_H (0x00000000)
value GRADIENT_FILL_RECT_V (0x00000001)
value GRADIENT_FILL_TRIANGLE (0x00000002)
value GRAY_BRUSH (2)
value GREEK_CHARSET (161)
value GROUP_NAME (0x80)
value GROUP_SECURITY_INFORMATION ((0x00000002L))
value GR_GDIOBJECTS (0)
value GR_GDIOBJECTS_PEAK (2)
value GR_GLOBAL (((HANDLE)-2))
value GR_USEROBJECTS (1)
value GR_USEROBJECTS_PEAK (4)
value GSS_ALLOW_INHERITED_COMMON (0x0001)
value GUID_CLASS_COMPORT (GUID_DEVINTERFACE_COMPORT)
value GUID_SERENUM_BUS_ENUMERATOR (GUID_DEVINTERFACE_SERENUM_BUS_ENUMERATOR)
value GUI_CARETBLINKING (0x00000001)
value GUI_INMENUMODE (0x00000004)
value GUI_INMOVESIZE (0x00000002)
value GUI_POPUPMENUMODE (0x00000010)
value GUI_SYSTEMMENUMODE (0x00000008)
value GWFS_INCLUDE_ANCESTORS (0x00000001)
value GWLP_HINSTANCE ((-6))
value GWLP_HWNDPARENT ((-8))
value GWLP_ID ((-12))
value GWLP_USERDATA ((-21))
value GWLP_WNDPROC ((-4))
value GWL_EXSTYLE ((-20))
value GWL_ID ((-12))
value GWL_STYLE ((-16))
value GW_CHILD (5)
value GW_ENABLEDPOPUP (6)
value GW_HWNDFIRST (0)
value GW_HWNDLAST (1)
value GW_HWNDNEXT (2)
value GW_HWNDPREV (3)
value GW_MAX (6)
value GW_OWNER (4)
value HALFTONE (4)
value HANDLE_FLAG_INHERIT (0x00000001)
value HANDLE_FLAG_PROTECT_FROM_CLOSE (0x00000002)
value HANGEUL_CHARSET (129)
value HANGUL_CHARSET (129)
value HANGUP_COMPLETE (0x05)
value HANGUP_PENDING (0x04)
value HBMMENU_CALLBACK (((HBITMAP) -1))
value HBMMENU_MBAR_CLOSE (((HBITMAP) 5))
value HBMMENU_MBAR_CLOSE_D (((HBITMAP) 6))
value HBMMENU_MBAR_MINIMIZE (((HBITMAP) 3))
value HBMMENU_MBAR_MINIMIZE_D (((HBITMAP) 7))
value HBMMENU_MBAR_RESTORE (((HBITMAP) 2))
value HBMMENU_POPUP_CLOSE (((HBITMAP) 8))
value HBMMENU_POPUP_MAXIMIZE (((HBITMAP) 10))
value HBMMENU_POPUP_MINIMIZE (((HBITMAP) 11))
value HBMMENU_POPUP_RESTORE (((HBITMAP) 9))
value HBMMENU_SYSTEM (((HBITMAP) 1))
value HCBT_ACTIVATE (5)
value HCBT_CLICKSKIPPED (6)
value HCBT_CREATEWND (3)
value HCBT_DESTROYWND (4)
value HCBT_KEYSKIPPED (7)
value HCBT_MINMAX (1)
value HCBT_MOVESIZE (0)
value HCBT_QS (2)
value HCBT_SETFOCUS (9)
value HCBT_SYSCOMMAND (8)
value HCCE_CURRENT_USER (((HCERTCHAINENGINE)NULL))
value HCCE_LOCAL_MACHINE (((HCERTCHAINENGINE)0x1))
value HCCE_SERIAL_LOCAL_MACHINE (((HCERTCHAINENGINE)0x2))
value HCF_AVAILABLE (0x00000002)
value HCF_CONFIRMHOTKEY (0x00000008)
value HCF_DEFAULTDESKTOP (0x00000200)
value HCF_HIGHCONTRASTON (0x00000001)
value HCF_HOTKEYACTIVE (0x00000004)
value HCF_HOTKEYAVAILABLE (0x00000040)
value HCF_HOTKEYSOUND (0x00000010)
value HCF_INDICATOR (0x00000020)
value HCF_LOGONDESKTOP (0x00000100)
value HCF_OPTION_NOTHEMECHANGE (0x00001000)
value HCN_E_ADAPTER_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0006L))
value HCN_E_ADDR_INVALID_OR_RESERVED (_HRESULT_TYPEDEF_(0x803B002FL))
value HCN_E_DEGRADED_OPERATION (_HRESULT_TYPEDEF_(0x803B0017L))
value HCN_E_ENDPOINT_ALREADY_ATTACHED (_HRESULT_TYPEDEF_(0x803B0014L))
value HCN_E_ENDPOINT_NAMESPACE_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x803B002BL))
value HCN_E_ENDPOINT_NOT_ATTACHED (_HRESULT_TYPEDEF_(0x803B0034L))
value HCN_E_ENDPOINT_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0002L))
value HCN_E_ENDPOINT_NOT_LOCAL (_HRESULT_TYPEDEF_(0x803B0035L))
value HCN_E_ENDPOINT_SHARING_DISABLED (_HRESULT_TYPEDEF_(0x803B001DL))
value HCN_E_ENTITY_HAS_REFERENCES (_HRESULT_TYPEDEF_(0x803B002CL))
value HCN_E_GUID_CONVERSION_FAILURE (_HRESULT_TYPEDEF_(0x803B0019L))
value HCN_E_ICS_DISABLED (_HRESULT_TYPEDEF_(0x803B002AL))
value HCN_E_INVALID_ENDPOINT (_HRESULT_TYPEDEF_(0x803B000CL))
value HCN_E_INVALID_INTERNAL_PORT (_HRESULT_TYPEDEF_(0x803B002DL))
value HCN_E_INVALID_IP (_HRESULT_TYPEDEF_(0x803B001EL))
value HCN_E_INVALID_IP_SUBNET (_HRESULT_TYPEDEF_(0x803B0033L))
value HCN_E_INVALID_JSON (_HRESULT_TYPEDEF_(0x803B001BL))
value HCN_E_INVALID_JSON_REFERENCE (_HRESULT_TYPEDEF_(0x803B001CL))
value HCN_E_INVALID_NETWORK (_HRESULT_TYPEDEF_(0x803B000AL))
value HCN_E_INVALID_NETWORK_TYPE (_HRESULT_TYPEDEF_(0x803B000BL))
value HCN_E_INVALID_POLICY (_HRESULT_TYPEDEF_(0x803B000DL))
value HCN_E_INVALID_POLICY_TYPE (_HRESULT_TYPEDEF_(0x803B000EL))
value HCN_E_INVALID_PREFIX (_HRESULT_TYPEDEF_(0x803B0030L))
value HCN_E_INVALID_REMOTE_ENDPOINT_OPERATION (_HRESULT_TYPEDEF_(0x803B000FL))
value HCN_E_INVALID_SUBNET (_HRESULT_TYPEDEF_(0x803B0032L))
value HCN_E_LAYER_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x803B0011L))
value HCN_E_LAYER_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0003L))
value HCN_E_MANAGER_STOPPED (_HRESULT_TYPEDEF_(0x803B0020L))
value HCN_E_MAPPING_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803B0016L))
value HCN_E_NAMESPACE_ATTACH_FAILED (_HRESULT_TYPEDEF_(0x803B002EL))
value HCN_E_NETWORK_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x803B0010L))
value HCN_E_NETWORK_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0001L))
value HCN_E_OBJECT_USED_AFTER_UNLOAD (_HRESULT_TYPEDEF_(0x803B0031L))
value HCN_E_POLICY_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x803B0012L))
value HCN_E_POLICY_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0008L))
value HCN_E_PORT_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x803B0013L))
value HCN_E_PORT_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0007L))
value HCN_E_REGKEY_FAILURE (_HRESULT_TYPEDEF_(0x803B001AL))
value HCN_E_REQUEST_UNSUPPORTED (_HRESULT_TYPEDEF_(0x803B0015L))
value HCN_E_SHARED_SWITCH_MODIFICATION (_HRESULT_TYPEDEF_(0x803B0018L))
value HCN_E_SUBNET_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0005L))
value HCN_E_SWITCH_EXTENSION_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B001FL))
value HCN_E_SWITCH_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0004L))
value HCN_E_VFP_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x803B0037L))
value HCN_E_VFP_PORTSETTING_NOT_FOUND (_HRESULT_TYPEDEF_(0x803B0009L))
value HCN_INTERFACEPARAMETERS_ALREADY_APPLIED (_HRESULT_TYPEDEF_(0x803B0036L))
value HCS_E_ACCESS_DENIED (_HRESULT_TYPEDEF_(0x8037011BL))
value HCS_E_CONNECTION_CLOSED (_HRESULT_TYPEDEF_(0x8037010AL))
value HCS_E_CONNECTION_TIMEOUT (_HRESULT_TYPEDEF_(0x80370109L))
value HCS_E_CONNECT_FAILED (_HRESULT_TYPEDEF_(0x80370108L))
value HCS_E_GUEST_CRITICAL_ERROR (_HRESULT_TYPEDEF_(0x8037011CL))
value HCS_E_HYPERV_NOT_INSTALLED (_HRESULT_TYPEDEF_(0x80370102L))
value HCS_E_IMAGE_MISMATCH (_HRESULT_TYPEDEF_(0x80370101L))
value HCS_E_INVALID_JSON (_HRESULT_TYPEDEF_(0x8037010DL))
value HCS_E_INVALID_LAYER (_HRESULT_TYPEDEF_(0x80370112L))
value HCS_E_INVALID_STATE (_HRESULT_TYPEDEF_(0x80370105L))
value HCS_E_OPERATION_ALREADY_CANCELLED (_HRESULT_TYPEDEF_(0x80370121L))
value HCS_E_OPERATION_ALREADY_STARTED (_HRESULT_TYPEDEF_(0x80370116L))
value HCS_E_OPERATION_NOT_STARTED (_HRESULT_TYPEDEF_(0x80370115L))
value HCS_E_OPERATION_PENDING (_HRESULT_TYPEDEF_(0x80370117L))
value HCS_E_OPERATION_RESULT_ALLOCATION_FAILED (_HRESULT_TYPEDEF_(0x8037011AL))
value HCS_E_OPERATION_SYSTEM_CALLBACK_ALREADY_SET (_HRESULT_TYPEDEF_(0x80370119L))
value HCS_E_OPERATION_TIMEOUT (_HRESULT_TYPEDEF_(0x80370118L))
value HCS_E_PROCESS_ALREADY_STOPPED (_HRESULT_TYPEDEF_(0x8037011FL))
value HCS_E_PROCESS_INFO_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x8037011DL))
value HCS_E_PROTOCOL_ERROR (_HRESULT_TYPEDEF_(0x80370111L))
value HCS_E_SERVICE_DISCONNECT (_HRESULT_TYPEDEF_(0x8037011EL))
value HCS_E_SERVICE_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x80370114L))
value HCS_E_SYSTEM_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x8037010FL))
value HCS_E_SYSTEM_ALREADY_STOPPED (_HRESULT_TYPEDEF_(0x80370110L))
value HCS_E_SYSTEM_NOT_CONFIGURED_FOR_OPERATION (_HRESULT_TYPEDEF_(0x80370120L))
value HCS_E_SYSTEM_NOT_FOUND (_HRESULT_TYPEDEF_(0x8037010EL))
value HCS_E_TERMINATED (_HRESULT_TYPEDEF_(0x80370107L))
value HCS_E_TERMINATED_DURING_START (_HRESULT_TYPEDEF_(0x80370100L))
value HCS_E_UNEXPECTED_EXIT (_HRESULT_TYPEDEF_(0x80370106L))
value HCS_E_UNKNOWN_MESSAGE (_HRESULT_TYPEDEF_(0x8037010BL))
value HCS_E_UNSUPPORTED_PROTOCOL_VERSION (_HRESULT_TYPEDEF_(0x8037010CL))
value HCS_E_WINDOWS_INSIDER_REQUIRED (_HRESULT_TYPEDEF_(0x80370113L))
value HC_ACTION (0)
value HC_GETNEXT (1)
value HC_NOREM (HC_NOREMOVE)
value HC_NOREMOVE (3)
value HC_SKIP (2)
value HC_SYSMODALOFF (5)
value HC_SYSMODALON (4)
value HDATA_APPOWNED (0x0001)
value HEAP_CREATE_ENABLE_EXECUTE (0x00040000)
value HEAP_CREATE_ENABLE_TRACING (0x00020000)
value HEAP_CREATE_HARDENED (0x00000200)
value HEAP_CREATE_SEGMENT_HEAP (0x00000100)
value HEAP_DISABLE_COALESCE_ON_FREE (0x00000080)
value HEAP_FREE_CHECKING_ENABLED (0x00000040)
value HEAP_GENERATE_EXCEPTIONS (0x00000004)
value HEAP_GROWABLE (0x00000002)
value HEAP_MAXIMUM_TAG (0x0FFF)
value HEAP_NO_SERIALIZE (0x00000001)
value HEAP_OPTIMIZE_RESOURCES_CURRENT_VERSION (1)
value HEAP_PSEUDO_TAG_FLAG (0x8000)
value HEAP_REALLOC_IN_PLACE_ONLY (0x00000010)
value HEAP_TAG_SHIFT (18)
value HEAP_TAIL_CHECKING_ENABLED (0x00000020)
value HEAP_ZERO_MEMORY (0x00000008)
value HEBREW_CHARSET (177)
value HELPINFO_MENUITEM (0x0002)
value HELPINFO_WINDOW (0x0001)
value HELPMSGSTRING (HELPMSGSTRINGA)
value HELP_COMMAND (0x0102L)
value HELP_CONTENTS (0x0003L)
value HELP_CONTEXT (0x0001L)
value HELP_CONTEXTMENU (0x000a)
value HELP_CONTEXTPOPUP (0x0008L)
value HELP_FINDER (0x000b)
value HELP_FORCEFILE (0x0009L)
value HELP_HELPONHELP (0x0004L)
value HELP_INDEX (0x0003L)
value HELP_KEY (0x0101L)
value HELP_MULTIKEY (0x0201L)
value HELP_PARTIALKEY (0x0105L)
value HELP_QUIT (0x0002L)
value HELP_SETCONTENTS (0x0005L)
value HELP_SETINDEX (0x0005L)
value HELP_SETPOPUP_POS (0x000d)
value HELP_SETWINPOS (0x0203L)
value HELP_TCARD (0x8000)
value HELP_TCARD_DATA (0x0010)
value HELP_TCARD_OTHER_CALLER (0x0011)
value HELP_WM_HELP (0x000c)
value HFILE_ERROR (((HFILE)-1))
value HIBERFILE_TYPE_FULL (0x02)
value HIBERFILE_TYPE_MAX (0x03)
value HIBERFILE_TYPE_NONE (0x00)
value HIBERFILE_TYPE_REDUCED (0x01)
value HIDE_WINDOW (0)
value HIGH_LEVEL (15)
value HIGH_PRIORITY_CLASS (0x00000080)
value HIGH_SURROGATE_END (0xdbff)
value HIGH_SURROGATE_START (0xd800)
value HINSTANCE_ERROR (32)
value HISTORY_NO_DUP_FLAG (0x1)
value HIST_NO_OF_BUCKETS (24)
value HKEY_CLASSES_ROOT ((( HKEY ) (ULONG_PTR)((LONG)0x80000000) ))
value HKEY_CURRENT_CONFIG ((( HKEY ) (ULONG_PTR)((LONG)0x80000005) ))
value HKEY_CURRENT_USER ((( HKEY ) (ULONG_PTR)((LONG)0x80000001) ))
value HKEY_CURRENT_USER_LOCAL_SETTINGS ((( HKEY ) (ULONG_PTR)((LONG)0x80000007) ))
value HKEY_DYN_DATA ((( HKEY ) (ULONG_PTR)((LONG)0x80000006) ))
value HKEY_LOCAL_MACHINE ((( HKEY ) (ULONG_PTR)((LONG)0x80000002) ))
value HKEY_PERFORMANCE_DATA ((( HKEY ) (ULONG_PTR)((LONG)0x80000004) ))
value HKEY_PERFORMANCE_NLSTEXT ((( HKEY ) (ULONG_PTR)((LONG)0x80000060) ))
value HKEY_PERFORMANCE_TEXT ((( HKEY ) (ULONG_PTR)((LONG)0x80000050) ))
value HKEY_USERS ((( HKEY ) (ULONG_PTR)((LONG)0x80000003) ))
value HKL_NEXT (1)
value HKL_PREV (0)
value HOLLOW_BRUSH (NULL_BRUSH)
value HORZRES (8)
value HORZSIZE (4)
value HOST_NOT_FOUND (WSAHOST_NOT_FOUND)
value HOVER_DEFAULT (0xFFFFFFFF)
value HP_ALGID (0x0001)
value HP_HASHSIZE (0x0004)
value HP_HASHVAL (0x0002)
value HP_HMAC_INFO (0x0005)
value HSHELL_ACCESSIBILITYSTATE (11)
value HSHELL_ACTIVATESHELLWINDOW (3)
value HSHELL_APPCOMMAND (12)
value HSHELL_ENDTASK (10)
value HSHELL_FLASH ((HSHELL_REDRAW|HSHELL_HIGHBIT))
value HSHELL_GETMINRECT (5)
value HSHELL_HIGHBIT (0x8000)
value HSHELL_LANGUAGE (8)
value HSHELL_MONITORCHANGED (16)
value HSHELL_REDRAW (6)
value HSHELL_RUDEAPPACTIVATED ((HSHELL_WINDOWACTIVATED|HSHELL_HIGHBIT))
value HSHELL_SYSMENU (9)
value HSHELL_TASKMAN (7)
value HSHELL_WINDOWACTIVATED (4)
value HSHELL_WINDOWCREATED (1)
value HSHELL_WINDOWDESTROYED (2)
value HSHELL_WINDOWREPLACED (13)
value HSHELL_WINDOWREPLACING (14)
value HSP_BASE_ERROR_MASK (_HRESULT_TYPEDEF_(0x81290100L))
value HSP_BASE_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x812901FFL))
value HSP_BS_ERROR_MASK (_HRESULT_TYPEDEF_(0x81281000L))
value HSP_BS_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x812810FFL))
value HSP_DRV_ERROR_MASK (_HRESULT_TYPEDEF_(0x81290000L))
value HSP_DRV_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x812900FFL))
value HSP_E_ERROR_MASK (_HRESULT_TYPEDEF_(0x81280000L))
value HSP_E_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x81280FFFL))
value HSP_KSP_ALGORITHM_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x81290209L))
value HSP_KSP_BUFFER_TOO_SMALL (_HRESULT_TYPEDEF_(0x81290205L))
value HSP_KSP_DEVICE_NOT_READY (_HRESULT_TYPEDEF_(0x81290201L))
value HSP_KSP_ERROR_MASK (_HRESULT_TYPEDEF_(0x81290200L))
value HSP_KSP_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x812902FFL))
value HSP_KSP_INVALID_DATA (_HRESULT_TYPEDEF_(0x81290207L))
value HSP_KSP_INVALID_FLAGS (_HRESULT_TYPEDEF_(0x81290208L))
value HSP_KSP_INVALID_KEY_HANDLE (_HRESULT_TYPEDEF_(0x81290203L))
value HSP_KSP_INVALID_KEY_TYPE (_HRESULT_TYPEDEF_(0x8129020CL))
value HSP_KSP_INVALID_PARAMETER (_HRESULT_TYPEDEF_(0x81290204L))
value HSP_KSP_INVALID_PROVIDER_HANDLE (_HRESULT_TYPEDEF_(0x81290202L))
value HSP_KSP_KEY_ALREADY_FINALIZED (_HRESULT_TYPEDEF_(0x8129020AL))
value HSP_KSP_KEY_EXISTS (_HRESULT_TYPEDEF_(0x81290215L))
value HSP_KSP_KEY_LOAD_FAIL (_HRESULT_TYPEDEF_(0x81290217L))
value HSP_KSP_KEY_MISSING (_HRESULT_TYPEDEF_(0x81290216L))
value HSP_KSP_KEY_NOT_FINALIZED (_HRESULT_TYPEDEF_(0x8129020BL))
value HSP_KSP_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x81290206L))
value HSP_KSP_NO_MEMORY (_HRESULT_TYPEDEF_(0x81290210L))
value HSP_KSP_NO_MORE_ITEMS (_HRESULT_TYPEDEF_(0x81290218L))
value HSP_KSP_PARAMETER_NOT_SET (_HRESULT_TYPEDEF_(0x81290211L))
value HS_API_MAX (12)
value HS_BDIAGONAL (3)
value HS_CROSS (4)
value HS_DIAGCROSS (5)
value HS_FDIAGONAL (2)
value HS_HORIZONTAL (0)
value HS_VERTICAL (1)
value HTBORDER (18)
value HTBOTTOM (15)
value HTBOTTOMLEFT (16)
value HTBOTTOMRIGHT (17)
value HTCAPTION (2)
value HTCLIENT (1)
value HTCLOSE (20)
value HTERROR ((-2))
value HTGROWBOX (4)
value HTHELP (21)
value HTHSCROLL (6)
value HTLEFT (10)
value HTMAXBUTTON (9)
value HTMENU (5)
value HTMINBUTTON (8)
value HTNOWHERE (0)
value HTOBJECT (19)
value HTREDUCE (HTMINBUTTON)
value HTRIGHT (11)
value HTSIZE (HTGROWBOX)
value HTSIZEFIRST (HTLEFT)
value HTSIZELAST (HTBOTTOMRIGHT)
value HTSYSMENU (3)
value HTTOP (12)
value HTTOPLEFT (13)
value HTTOPRIGHT (14)
value HTTP_E_STATUS_AMBIGUOUS (_HRESULT_TYPEDEF_(0x8019012CL))
value HTTP_E_STATUS_BAD_GATEWAY (_HRESULT_TYPEDEF_(0x801901F6L))
value HTTP_E_STATUS_BAD_METHOD (_HRESULT_TYPEDEF_(0x80190195L))
value HTTP_E_STATUS_BAD_REQUEST (_HRESULT_TYPEDEF_(0x80190190L))
value HTTP_E_STATUS_CONFLICT (_HRESULT_TYPEDEF_(0x80190199L))
value HTTP_E_STATUS_DENIED (_HRESULT_TYPEDEF_(0x80190191L))
value HTTP_E_STATUS_EXPECTATION_FAILED (_HRESULT_TYPEDEF_(0x801901A1L))
value HTTP_E_STATUS_FORBIDDEN (_HRESULT_TYPEDEF_(0x80190193L))
value HTTP_E_STATUS_GATEWAY_TIMEOUT (_HRESULT_TYPEDEF_(0x801901F8L))
value HTTP_E_STATUS_GONE (_HRESULT_TYPEDEF_(0x8019019AL))
value HTTP_E_STATUS_LENGTH_REQUIRED (_HRESULT_TYPEDEF_(0x8019019BL))
value HTTP_E_STATUS_MOVED (_HRESULT_TYPEDEF_(0x8019012DL))
value HTTP_E_STATUS_NONE_ACCEPTABLE (_HRESULT_TYPEDEF_(0x80190196L))
value HTTP_E_STATUS_NOT_FOUND (_HRESULT_TYPEDEF_(0x80190194L))
value HTTP_E_STATUS_NOT_MODIFIED (_HRESULT_TYPEDEF_(0x80190130L))
value HTTP_E_STATUS_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x801901F5L))
value HTTP_E_STATUS_PAYMENT_REQ (_HRESULT_TYPEDEF_(0x80190192L))
value HTTP_E_STATUS_PRECOND_FAILED (_HRESULT_TYPEDEF_(0x8019019CL))
value HTTP_E_STATUS_PROXY_AUTH_REQ (_HRESULT_TYPEDEF_(0x80190197L))
value HTTP_E_STATUS_RANGE_NOT_SATISFIABLE (_HRESULT_TYPEDEF_(0x801901A0L))
value HTTP_E_STATUS_REDIRECT (_HRESULT_TYPEDEF_(0x8019012EL))
value HTTP_E_STATUS_REDIRECT_KEEP_VERB (_HRESULT_TYPEDEF_(0x80190133L))
value HTTP_E_STATUS_REDIRECT_METHOD (_HRESULT_TYPEDEF_(0x8019012FL))
value HTTP_E_STATUS_REQUEST_TIMEOUT (_HRESULT_TYPEDEF_(0x80190198L))
value HTTP_E_STATUS_REQUEST_TOO_LARGE (_HRESULT_TYPEDEF_(0x8019019DL))
value HTTP_E_STATUS_SERVER_ERROR (_HRESULT_TYPEDEF_(0x801901F4L))
value HTTP_E_STATUS_SERVICE_UNAVAIL (_HRESULT_TYPEDEF_(0x801901F7L))
value HTTP_E_STATUS_UNEXPECTED (_HRESULT_TYPEDEF_(0x80190001L))
value HTTP_E_STATUS_UNEXPECTED_CLIENT_ERROR (_HRESULT_TYPEDEF_(0x80190004L))
value HTTP_E_STATUS_UNEXPECTED_REDIRECTION (_HRESULT_TYPEDEF_(0x80190003L))
value HTTP_E_STATUS_UNEXPECTED_SERVER_ERROR (_HRESULT_TYPEDEF_(0x80190005L))
value HTTP_E_STATUS_UNSUPPORTED_MEDIA (_HRESULT_TYPEDEF_(0x8019019FL))
value HTTP_E_STATUS_URI_TOO_LONG (_HRESULT_TYPEDEF_(0x8019019EL))
value HTTP_E_STATUS_USE_PROXY (_HRESULT_TYPEDEF_(0x80190131L))
value HTTP_E_STATUS_VERSION_NOT_SUP (_HRESULT_TYPEDEF_(0x801901F9L))
value HTTRANSPARENT ((-1))
value HTVSCROLL (7)
value HTZOOM (HTMAXBUTTON)
value HWND_BOTTOM (((HWND)1))
value HWND_DESKTOP (((HWND)0))
value HWND_MESSAGE (((HWND)-3))
value HWND_NOTOPMOST (((HWND)-2))
value HWND_TOP (((HWND)0))
value HWND_TOPMOST (((HWND)-1))
value HW_PROFILE_GUIDLEN (39)
value IACE_CHILDREN (0x0001)
value IACE_DEFAULT (0x0010)
value IACE_IGNORENOCONTEXT (0x0020)
value ICMENUMPROC (ICMENUMPROCA)
value ICM_ADDPROFILE (1)
value ICM_DELETEPROFILE (2)
value ICM_DONE_OUTSIDEDC (4)
value ICM_OFF (1)
value ICM_ON (2)
value ICM_QUERY (3)
value ICM_QUERYMATCH (7)
value ICM_QUERYPROFILE (3)
value ICM_REGISTERICMATCHER (5)
value ICM_SETDEFAULTPROFILE (4)
value ICM_UNREGISTERICMATCHER (6)
value ICON_BIG (1)
value ICON_SMALL (0)
value IDABORT (3)
value IDANI_CAPTION (3)
value IDANI_OPEN (1)
value IDCANCEL (2)
value IDCLOSE (8)
value IDCONTINUE (11)
value IDC_APPSTARTING (MAKEINTRESOURCE(32650))
value IDC_ARROW (MAKEINTRESOURCE(32512))
value IDC_CROSS (MAKEINTRESOURCE(32515))
value IDC_HAND (MAKEINTRESOURCE(32649))
value IDC_HELP (MAKEINTRESOURCE(32651))
value IDC_IBEAM (MAKEINTRESOURCE(32513))
value IDC_ICON (MAKEINTRESOURCE(32641))
value IDC_MANAGE_LINK (1592)
value IDC_NO (MAKEINTRESOURCE(32648))
value IDC_PERSON (MAKEINTRESOURCE(32672))
value IDC_PIN (MAKEINTRESOURCE(32671))
value IDC_SIZE (MAKEINTRESOURCE(32640))
value IDC_SIZEALL (MAKEINTRESOURCE(32646))
value IDC_SIZENESW (MAKEINTRESOURCE(32643))
value IDC_SIZENS (MAKEINTRESOURCE(32645))
value IDC_SIZENWSE (MAKEINTRESOURCE(32642))
value IDC_SIZEWE (MAKEINTRESOURCE(32644))
value IDC_UPARROW (MAKEINTRESOURCE(32516))
value IDC_WAIT (MAKEINTRESOURCE(32514))
value IDENTIFY_BUFFER_SIZE (512)
value IDHELP (9)
value IDHOT_SNAPDESKTOP ((-2))
value IDHOT_SNAPWINDOW ((-1))
value IDH_CANCEL (28444)
value IDH_GENERIC_HELP_BUTTON (28442)
value IDH_HELP (28445)
value IDH_MISSING_CONTEXT (28441)
value IDH_NO_HELP (28440)
value IDH_OK (28443)
value IDIGNORE (5)
value IDI_APPLICATION (MAKEINTRESOURCE(32512))
value IDI_ASTERISK (MAKEINTRESOURCE(32516))
value IDI_ERROR (IDI_HAND)
value IDI_EXCLAMATION (MAKEINTRESOURCE(32515))
value IDI_HAND (MAKEINTRESOURCE(32513))
value IDI_INFORMATION (IDI_ASTERISK)
value IDI_QUESTION (MAKEINTRESOURCE(32514))
value IDI_SHIELD (MAKEINTRESOURCE(32518))
value IDI_WARNING (IDI_EXCLAMATION)
value IDI_WINLOGO (MAKEINTRESOURCE(32517))
value IDLE_PRIORITY_CLASS (0x00000040)
value IDLFLAG_FIN (( PARAMFLAG_FIN ))
value IDLFLAG_FLCID (( PARAMFLAG_FLCID ))
value IDLFLAG_FOUT (( PARAMFLAG_FOUT ))
value IDLFLAG_FRETVAL (( PARAMFLAG_FRETVAL ))
value IDLFLAG_NONE (( PARAMFLAG_NONE ))
value IDNO (7)
value IDN_ALLOW_UNASSIGNED (0x01)
value IDN_EMAIL_ADDRESS (0x04)
value IDN_RAW_PUNYCODE (0x08)
value IDOK (1)
value IDRETRY (4)
value IDTIMEOUT (32000)
value IDTRYAGAIN (10)
value IDYES (6)
value ID_CMD (0xEC)
value ID_DEFAULTINST (-2)
value ID_PSREBOOTSYSTEM ((ID_PSRESTARTWINDOWS | 0x1))
value ID_PSRESTARTWINDOWS (0x2)
value IE_BADID ((-1))
value IE_BAUDRATE ((-12))
value IE_BYTESIZE ((-11))
value IE_DEFAULT ((-5))
value IE_HARDWARE ((-10))
value IE_MEMORY ((-4))
value IE_NOPEN ((-3))
value IE_OPEN ((-2))
value IFX_RSA_KEYGEN_VUL_NOT_AFFECTED (0)
value IGIMIF_RIGHTMENU (0x0001)
value IGIMII_CMODE (0x0001)
value IGIMII_CONFIGURE (0x0004)
value IGIMII_HELP (0x0010)
value IGIMII_INPUTTOOLS (0x0040)
value IGIMII_OTHER (0x0020)
value IGIMII_SMODE (0x0002)
value IGIMII_TOOLS (0x0008)
value IGNORE (0)
value IGP_CONVERSION (0x00000008)
value IGP_GETIMEVERSION ((DWORD)(-4))
value IGP_PROPERTY (0x00000004)
value IGP_SELECT (0x00000018)
value IGP_SENTENCE (0x0000000c)
value IGP_SETCOMPSTR (0x00000014)
value IGP_UI (0x00000010)
value IID_NULL (GUID_NULL)
value ILLUMINANT_A (1)
value ILLUMINANT_B (2)
value ILLUMINANT_C (3)
value ILLUMINANT_DAYLIGHT (ILLUMINANT_C)
value ILLUMINANT_DEVICE_DEFAULT (0)
value ILLUMINANT_FLUORESCENT (ILLUMINANT_F2)
value ILLUMINANT_MAX_INDEX (ILLUMINANT_F2)
value ILLUMINANT_NTSC (ILLUMINANT_C)
value ILLUMINANT_TUNGSTEN (ILLUMINANT_A)
value IMAGE_ARCHIVE_START_SIZE (8)
value IMAGE_BITMAP (0)
value IMAGE_COMDAT_SELECT_ANY (2)
value IMAGE_COMDAT_SELECT_ASSOCIATIVE (5)
value IMAGE_COMDAT_SELECT_EXACT_MATCH (4)
value IMAGE_COMDAT_SELECT_LARGEST (6)
value IMAGE_COMDAT_SELECT_NEWEST (7)
value IMAGE_COMDAT_SELECT_NODUPLICATES (1)
value IMAGE_COMDAT_SELECT_SAME_SIZE (3)
value IMAGE_CURSOR (2)
value IMAGE_DEBUG_MISC_EXENAME (1)
value IMAGE_DEBUG_TYPE_BBT (IMAGE_DEBUG_TYPE_RESERVED10)
value IMAGE_DEBUG_TYPE_BORLAND (9)
value IMAGE_DEBUG_TYPE_CLSID (11)
value IMAGE_DEBUG_TYPE_CODEVIEW (2)
value IMAGE_DEBUG_TYPE_COFF (1)
value IMAGE_DEBUG_TYPE_EXCEPTION (5)
value IMAGE_DEBUG_TYPE_EX_DLLCHARACTERISTICS (20)
value IMAGE_DEBUG_TYPE_FIXUP (6)
value IMAGE_DEBUG_TYPE_FPO (3)
value IMAGE_DEBUG_TYPE_ILTCG (14)
value IMAGE_DEBUG_TYPE_MISC (4)
value IMAGE_DEBUG_TYPE_MPX (15)
value IMAGE_DEBUG_TYPE_OMAP_FROM_SRC (8)
value IMAGE_DEBUG_TYPE_OMAP_TO_SRC (7)
value IMAGE_DEBUG_TYPE_POGO (13)
value IMAGE_DEBUG_TYPE_REPRO (16)
value IMAGE_DEBUG_TYPE_SPGO (18)
value IMAGE_DEBUG_TYPE_UNKNOWN (0)
value IMAGE_DEBUG_TYPE_VC_FEATURE (12)
value IMAGE_DIRECTORY_ENTRY_ARCHITECTURE (7)
value IMAGE_DIRECTORY_ENTRY_BASERELOC (5)
value IMAGE_DIRECTORY_ENTRY_BOUND_IMPORT (11)
value IMAGE_DIRECTORY_ENTRY_COM_DESCRIPTOR (14)
value IMAGE_DIRECTORY_ENTRY_DEBUG (6)
value IMAGE_DIRECTORY_ENTRY_DELAY_IMPORT (13)
value IMAGE_DIRECTORY_ENTRY_EXCEPTION (3)
value IMAGE_DIRECTORY_ENTRY_EXPORT (0)
value IMAGE_DIRECTORY_ENTRY_GLOBALPTR (8)
value IMAGE_DIRECTORY_ENTRY_IAT (12)
value IMAGE_DIRECTORY_ENTRY_IMPORT (1)
value IMAGE_DIRECTORY_ENTRY_LOAD_CONFIG (10)
value IMAGE_DIRECTORY_ENTRY_RESOURCE (2)
value IMAGE_DIRECTORY_ENTRY_SECURITY (4)
value IMAGE_DIRECTORY_ENTRY_TLS (9)
value IMAGE_DLLCHARACTERISTICS_APPCONTAINER (0x1000)
value IMAGE_DLLCHARACTERISTICS_DYNAMIC_BASE (0x0040)
value IMAGE_DLLCHARACTERISTICS_EX_CET_COMPAT (0x01)
value IMAGE_DLLCHARACTERISTICS_EX_CET_COMPAT_STRICT_MODE (0x02)
value IMAGE_DLLCHARACTERISTICS_EX_CET_DYNAMIC_APIS_ALLOW_IN_PROC (0x08)
value IMAGE_DLLCHARACTERISTICS_EX_CET_SET_CONTEXT_IP_VALIDATION_RELAXED_MODE (0x04)
value IMAGE_DLLCHARACTERISTICS_FORCE_INTEGRITY (0x0080)
value IMAGE_DLLCHARACTERISTICS_GUARD_CF (0x4000)
value IMAGE_DLLCHARACTERISTICS_HIGH_ENTROPY_VA (0x0020)
value IMAGE_DLLCHARACTERISTICS_NO_BIND (0x0800)
value IMAGE_DLLCHARACTERISTICS_NO_ISOLATION (0x0200)
value IMAGE_DLLCHARACTERISTICS_NO_SEH (0x0400)
value IMAGE_DLLCHARACTERISTICS_NX_COMPAT (0x0100)
value IMAGE_DLLCHARACTERISTICS_TERMINAL_SERVER_AWARE (0x8000)
value IMAGE_DLLCHARACTERISTICS_WDM_DRIVER (0x2000)
value IMAGE_DOS_SIGNATURE (0x5A4D)
value IMAGE_DYNAMIC_RELOCATION_FUNCTION_OVERRIDE (0x00000007)
value IMAGE_DYNAMIC_RELOCATION_GUARD_IMPORT_CONTROL_TRANSFER (0x00000003)
value IMAGE_DYNAMIC_RELOCATION_GUARD_INDIR_CONTROL_TRANSFER (0x00000004)
value IMAGE_DYNAMIC_RELOCATION_GUARD_RF_EPILOGUE (0x00000002)
value IMAGE_DYNAMIC_RELOCATION_GUARD_RF_PROLOGUE (0x00000001)
value IMAGE_DYNAMIC_RELOCATION_GUARD_SWITCHTABLE_BRANCH (0x00000005)
value IMAGE_ENCLAVE_FLAG_PRIMARY_IMAGE (0x00000001)
value IMAGE_ENCLAVE_IMPORT_MATCH_AUTHOR_ID (0x00000002)
value IMAGE_ENCLAVE_IMPORT_MATCH_FAMILY_ID (0x00000003)
value IMAGE_ENCLAVE_IMPORT_MATCH_IMAGE_ID (0x00000004)
value IMAGE_ENCLAVE_IMPORT_MATCH_NONE (0x00000000)
value IMAGE_ENCLAVE_IMPORT_MATCH_UNIQUE_ID (0x00000001)
value IMAGE_ENCLAVE_LONG_ID_LENGTH (ENCLAVE_LONG_ID_LENGTH)
value IMAGE_ENCLAVE_POLICY_DEBUGGABLE (0x00000001)
value IMAGE_ENCLAVE_SHORT_ID_LENGTH (ENCLAVE_SHORT_ID_LENGTH)
value IMAGE_ENHMETAFILE (3)
value IMAGE_FILE_AGGRESIVE_WS_TRIM (0x0010)
value IMAGE_FILE_BYTES_REVERSED_HI (0x8000)
value IMAGE_FILE_BYTES_REVERSED_LO (0x0080)
value IMAGE_FILE_DEBUG_STRIPPED (0x0200)
value IMAGE_FILE_DLL (0x2000)
value IMAGE_FILE_EXECUTABLE_IMAGE (0x0002)
value IMAGE_FILE_LARGE_ADDRESS_AWARE (0x0020)
value IMAGE_FILE_LINE_NUMS_STRIPPED (0x0004)
value IMAGE_FILE_LOCAL_SYMS_STRIPPED (0x0008)
value IMAGE_FILE_MACHINE_ALPHA (0x0184)
value IMAGE_FILE_MACHINE_ARM (0x01c0)
value IMAGE_FILE_MACHINE_ARMNT (0x01c4)
value IMAGE_FILE_MACHINE_CEE (0xC0EE)
value IMAGE_FILE_MACHINE_CEF (0x0CEF)
value IMAGE_FILE_MACHINE_EBC (0x0EBC)
value IMAGE_FILE_MACHINE_MIPSFPU (0x0366)
value IMAGE_FILE_MACHINE_POWERPC (0x01F0)
value IMAGE_FILE_MACHINE_POWERPCFP (0x01f1)
value IMAGE_FILE_MACHINE_TARGET_HOST (0x0001)
value IMAGE_FILE_MACHINE_THUMB (0x01c2)
value IMAGE_FILE_MACHINE_TRICORE (0x0520)
value IMAGE_FILE_MACHINE_UNKNOWN (0)
value IMAGE_FILE_NET_RUN_FROM_SWAP (0x0800)
value IMAGE_FILE_RELOCS_STRIPPED (0x0001)
value IMAGE_FILE_REMOVABLE_RUN_FROM_SWAP (0x0400)
value IMAGE_FILE_SYSTEM (0x1000)
value IMAGE_FILE_UP_SYSTEM_ONLY (0x4000)
value IMAGE_FUNCTION_OVERRIDE_INVALID (0)
value IMAGE_GUARD_CASTGUARD_PRESENT (0x01000000)
value IMAGE_GUARD_CFW_INSTRUMENTED (0x00000200)
value IMAGE_GUARD_CF_ENABLE_EXPORT_SUPPRESSION (0x00008000)
value IMAGE_GUARD_CF_EXPORT_SUPPRESSION_INFO_PRESENT (0x00004000)
value IMAGE_GUARD_CF_FUNCTION_TABLE_PRESENT (0x00000400)
value IMAGE_GUARD_CF_FUNCTION_TABLE_SIZE_MASK (0xF0000000)
value IMAGE_GUARD_CF_FUNCTION_TABLE_SIZE_SHIFT (28)
value IMAGE_GUARD_CF_INSTRUMENTED (0x00000100)
value IMAGE_GUARD_CF_LONGJUMP_TABLE_PRESENT (0x00010000)
value IMAGE_GUARD_DELAYLOAD_IAT_IN_ITS_OWN_SECTION (0x00002000)
value IMAGE_GUARD_EH_CONTINUATION_TABLE_PRESENT (0x00400000)
value IMAGE_GUARD_FLAG_EXPORT_SUPPRESSED (0x02)
value IMAGE_GUARD_FLAG_FID_LANGEXCPTHANDLER (0x04)
value IMAGE_GUARD_FLAG_FID_SUPPRESSED (0x01)
value IMAGE_GUARD_FLAG_FID_XFG (0x08)
value IMAGE_GUARD_MEMCPY_PRESENT (0x02000000)
value IMAGE_GUARD_PROTECT_DELAYLOAD_IAT (0x00001000)
value IMAGE_GUARD_RETPOLINE_PRESENT (0x00100000)
value IMAGE_GUARD_RF_ENABLE (0x00040000)
value IMAGE_GUARD_RF_INSTRUMENTED (0x00020000)
value IMAGE_GUARD_RF_STRICT (0x00080000)
value IMAGE_GUARD_SECURITY_COOKIE_UNUSED (0x00000800)
value IMAGE_GUARD_XFG_ENABLED (0x00800000)
value IMAGE_HOT_PATCH_ABSOLUTE (0x0002C000)
value IMAGE_HOT_PATCH_BASE_CAN_ROLL_BACK (0x00000002)
value IMAGE_HOT_PATCH_BASE_OBLIGATORY (0x00000001)
value IMAGE_HOT_PATCH_CALL_TARGET (0x00044000)
value IMAGE_HOT_PATCH_CHUNK_INVERSE (0x80000000)
value IMAGE_HOT_PATCH_CHUNK_OBLIGATORY (0x40000000)
value IMAGE_HOT_PATCH_CHUNK_RESERVED (0x3FF03000)
value IMAGE_HOT_PATCH_CHUNK_SIZE (0x00000FFF)
value IMAGE_HOT_PATCH_CHUNK_SOURCE_RVA (0x00008000)
value IMAGE_HOT_PATCH_CHUNK_TARGET_RVA (0x00004000)
value IMAGE_HOT_PATCH_CHUNK_TYPE (0x000FC000)
value IMAGE_HOT_PATCH_DYNAMIC_VALUE (0x00078000)
value IMAGE_HOT_PATCH_FUNCTION (0x0001C000)
value IMAGE_HOT_PATCH_INDIRECT (0x0005C000)
value IMAGE_HOT_PATCH_NONE (0x00000000)
value IMAGE_HOT_PATCH_NO_CALL_TARGET (0x00064000)
value IMAGE_ICON (1)
value IMAGE_NT_OPTIONAL_HDR_MAGIC (IMAGE_NT_OPTIONAL_HDR64_MAGIC)
value IMAGE_NT_SIGNATURE (0x00004550)
value IMAGE_NUMBEROF_DIRECTORY_ENTRIES (16)
value IMAGE_ORDINAL_FLAG (IMAGE_ORDINAL_FLAG64)
value IMAGE_POLICY_METADATA_VERSION (1)
value IMAGE_REL_ALPHA_ABSOLUTE (0x0000)
value IMAGE_REL_ALPHA_BRADDR (0x0007)
value IMAGE_REL_ALPHA_GPDISP (0x0006)
value IMAGE_REL_ALPHA_GPRELHI (0x0017)
value IMAGE_REL_ALPHA_GPRELLO (0x0016)
value IMAGE_REL_ALPHA_HINT (0x0008)
value IMAGE_REL_ALPHA_INLINE_REFLONG (0x0009)
value IMAGE_REL_ALPHA_LITERAL (0x0004)
value IMAGE_REL_ALPHA_LITUSE (0x0005)
value IMAGE_REL_ALPHA_MATCH (0x000D)
value IMAGE_REL_ALPHA_PAIR (0x000C)
value IMAGE_REL_ALPHA_REFHI (0x000A)
value IMAGE_REL_ALPHA_REFLO (0x000B)
value IMAGE_REL_ALPHA_REFLONG (0x0001)
value IMAGE_REL_ALPHA_REFLONGNB (0x0010)
value IMAGE_REL_ALPHA_REFQUAD (0x0002)
value IMAGE_REL_ALPHA_SECREL (0x000F)
value IMAGE_REL_ALPHA_SECRELHI (0x0012)
value IMAGE_REL_ALPHA_SECRELLO (0x0011)
value IMAGE_REL_ALPHA_SECTION (0x000E)
value IMAGE_REL_AM_ABSOLUTE (0x0000)
value IMAGE_REL_AM_FUNCINFO (0x0004)
value IMAGE_REL_AM_SECREL (0x0007)
value IMAGE_REL_AM_SECTION (0x0008)
value IMAGE_REL_AM_TOKEN (0x0009)
value IMAGE_REL_ARM_ABSOLUTE (0x0000)
value IMAGE_REL_ARM_SECREL (0x000F)
value IMAGE_REL_ARM_SECTION (0x000E)
value IMAGE_REL_ARM_TOKEN (0x0005)
value IMAGE_REL_BASED_ABSOLUTE (0)
value IMAGE_REL_BASED_HIGH (1)
value IMAGE_REL_BASED_HIGHADJ (4)
value IMAGE_REL_BASED_HIGHLOW (3)
value IMAGE_REL_BASED_LOW (2)
value IMAGE_REL_BASED_MIPS_JMPADDR (5)
value IMAGE_REL_BASED_RESERVED (6)
value IMAGE_REL_CEE_ABSOLUTE (0x0000)
value IMAGE_REL_CEE_SECREL (0x0005)
value IMAGE_REL_CEE_SECTION (0x0004)
value IMAGE_REL_CEE_TOKEN (0x0006)
value IMAGE_REL_CEF_ABSOLUTE (0x0000)
value IMAGE_REL_CEF_SECREL (0x0005)
value IMAGE_REL_CEF_SECTION (0x0004)
value IMAGE_REL_CEF_TOKEN (0x0006)
value IMAGE_REL_EBC_ABSOLUTE (0x0000)
value IMAGE_REL_EBC_SECREL (0x0004)
value IMAGE_REL_EBC_SECTION (0x0003)
value IMAGE_REL_MIPS_ABSOLUTE (0x0000)
value IMAGE_REL_MIPS_GPREL (0x0006)
value IMAGE_REL_MIPS_JMPADDR (0x0003)
value IMAGE_REL_MIPS_LITERAL (0x0007)
value IMAGE_REL_MIPS_PAIR (0x0025)
value IMAGE_REL_MIPS_REFHALF (0x0001)
value IMAGE_REL_MIPS_REFHI (0x0004)
value IMAGE_REL_MIPS_REFLO (0x0005)
value IMAGE_REL_MIPS_REFWORD (0x0002)
value IMAGE_REL_MIPS_REFWORDNB (0x0022)
value IMAGE_REL_MIPS_SECREL (0x000B)
value IMAGE_REL_MIPS_SECRELHI (0x000D)
value IMAGE_REL_MIPS_SECRELLO (0x000C)
value IMAGE_REL_MIPS_SECTION (0x000A)
value IMAGE_REL_MIPS_TOKEN (0x000E)
value IMAGE_REL_PPC_ABSOLUTE (0x0000)
value IMAGE_REL_PPC_BRNTAKEN (0x0400)
value IMAGE_REL_PPC_BRTAKEN (0x0200)
value IMAGE_REL_PPC_GPREL (0x0015)
value IMAGE_REL_PPC_IFGLUE (0x000D)
value IMAGE_REL_PPC_IMGLUE (0x000E)
value IMAGE_REL_PPC_NEG (0x0100)
value IMAGE_REL_PPC_PAIR (0x0012)
value IMAGE_REL_PPC_REFHI (0x0010)
value IMAGE_REL_PPC_REFLO (0x0011)
value IMAGE_REL_PPC_SECREL (0x000B)
value IMAGE_REL_PPC_SECRELHI (0x0014)
value IMAGE_REL_PPC_SECRELLO (0x0013)
value IMAGE_REL_PPC_SECTION (0x000C)
value IMAGE_REL_PPC_TOCDEFN (0x0800)
value IMAGE_REL_PPC_TOKEN (0x0016)
value IMAGE_REL_PPC_TYPEMASK (0x00FF)
value IMAGE_REL_SHM_PAIR (0x0018)
value IMAGE_REL_SHM_PCRELPT (0x0013)
value IMAGE_REL_SHM_REFHALF (0x0015)
value IMAGE_REL_SHM_REFLO (0x0014)
value IMAGE_REL_SHM_RELHALF (0x0017)
value IMAGE_REL_SHM_RELLO (0x0016)
value IMAGE_REL_SH_NOMODE (0x8000)
value IMAGE_RESOURCE_DATA_IS_DIRECTORY (0x80000000)
value IMAGE_RESOURCE_NAME_IS_STRING (0x80000000)
value IMAGE_ROM_OPTIONAL_HDR_MAGIC (0x107)
value IMAGE_SCN_ALIGN_MASK (0x00F00000)
value IMAGE_SCN_CNT_CODE (0x00000020)
value IMAGE_SCN_CNT_INITIALIZED_DATA (0x00000040)
value IMAGE_SCN_CNT_UNINITIALIZED_DATA (0x00000080)
value IMAGE_SCN_GPREL (0x00008000)
value IMAGE_SCN_LNK_COMDAT (0x00001000)
value IMAGE_SCN_LNK_INFO (0x00000200)
value IMAGE_SCN_LNK_NRELOC_OVFL (0x01000000)
value IMAGE_SCN_LNK_OTHER (0x00000100)
value IMAGE_SCN_LNK_REMOVE (0x00000800)
value IMAGE_SCN_MEM_DISCARDABLE (0x02000000)
value IMAGE_SCN_MEM_EXECUTE (0x20000000)
value IMAGE_SCN_MEM_FARDATA (0x00008000)
value IMAGE_SCN_MEM_LOCKED (0x00040000)
value IMAGE_SCN_MEM_NOT_CACHED (0x04000000)
value IMAGE_SCN_MEM_NOT_PAGED (0x08000000)
value IMAGE_SCN_MEM_PRELOAD (0x00080000)
value IMAGE_SCN_MEM_PURGEABLE (0x00020000)
value IMAGE_SCN_MEM_READ (0x40000000)
value IMAGE_SCN_MEM_SHARED (0x10000000)
value IMAGE_SCN_MEM_WRITE (0x80000000)
value IMAGE_SCN_NO_DEFER_SPEC_EXC (0x00004000)
value IMAGE_SCN_SCALE_INDEX (0x00000001)
value IMAGE_SCN_TYPE_NO_PAD (0x00000008)
value IMAGE_SEPARATE_DEBUG_FLAGS_MASK (0x8000)
value IMAGE_SEPARATE_DEBUG_MISMATCH (0x8000)
value IMAGE_SEPARATE_DEBUG_SIGNATURE (0x4944)
value IMAGE_SIZEOF_ARCHIVE_MEMBER_HDR (60)
value IMAGE_SIZEOF_FILE_HEADER (20)
value IMAGE_SIZEOF_SECTION_HEADER (40)
value IMAGE_SIZEOF_SHORT_NAME (8)
value IMAGE_SIZEOF_SYMBOL (18)
value IMAGE_SUBSYSTEM_EFI_APPLICATION (10)
value IMAGE_SUBSYSTEM_EFI_BOOT_SERVICE_DRIVER (11)
value IMAGE_SUBSYSTEM_EFI_ROM (13)
value IMAGE_SUBSYSTEM_EFI_RUNTIME_DRIVER (12)
value IMAGE_SUBSYSTEM_NATIVE (1)
value IMAGE_SUBSYSTEM_NATIVE_WINDOWS (8)
value IMAGE_SUBSYSTEM_POSIX_CUI (7)
value IMAGE_SUBSYSTEM_UNKNOWN (0)
value IMAGE_SUBSYSTEM_WINDOWS_BOOT_APPLICATION (16)
value IMAGE_SUBSYSTEM_WINDOWS_CE_GUI (9)
value IMAGE_SUBSYSTEM_WINDOWS_CUI (3)
value IMAGE_SUBSYSTEM_WINDOWS_GUI (2)
value IMAGE_SUBSYSTEM_XBOX (14)
value IMAGE_SUBSYSTEM_XBOX_CODE_CATALOG (17)
value IMAGE_SYM_ABSOLUTE ((SHORT)-1)
value IMAGE_SYM_CLASS_ARGUMENT (0x0009)
value IMAGE_SYM_CLASS_AUTOMATIC (0x0001)
value IMAGE_SYM_CLASS_BIT_FIELD (0x0012)
value IMAGE_SYM_CLASS_BLOCK (0x0064)
value IMAGE_SYM_CLASS_CLR_TOKEN (0x006B)
value IMAGE_SYM_CLASS_END_OF_FUNCTION ((BYTE )-1)
value IMAGE_SYM_CLASS_END_OF_STRUCT (0x0066)
value IMAGE_SYM_CLASS_ENUM_TAG (0x000F)
value IMAGE_SYM_CLASS_EXTERNAL (0x0002)
value IMAGE_SYM_CLASS_EXTERNAL_DEF (0x0005)
value IMAGE_SYM_CLASS_FAR_EXTERNAL (0x0044)
value IMAGE_SYM_CLASS_FILE (0x0067)
value IMAGE_SYM_CLASS_FUNCTION (0x0065)
value IMAGE_SYM_CLASS_LABEL (0x0006)
value IMAGE_SYM_CLASS_MEMBER_OF_ENUM (0x0010)
value IMAGE_SYM_CLASS_MEMBER_OF_STRUCT (0x0008)
value IMAGE_SYM_CLASS_MEMBER_OF_UNION (0x000B)
value IMAGE_SYM_CLASS_NULL (0x0000)
value IMAGE_SYM_CLASS_REGISTER (0x0004)
value IMAGE_SYM_CLASS_REGISTER_PARAM (0x0011)
value IMAGE_SYM_CLASS_SECTION (0x0068)
value IMAGE_SYM_CLASS_STATIC (0x0003)
value IMAGE_SYM_CLASS_STRUCT_TAG (0x000A)
value IMAGE_SYM_CLASS_TYPE_DEFINITION (0x000D)
value IMAGE_SYM_CLASS_UNDEFINED_LABEL (0x0007)
value IMAGE_SYM_CLASS_UNDEFINED_STATIC (0x000E)
value IMAGE_SYM_CLASS_UNION_TAG (0x000C)
value IMAGE_SYM_CLASS_WEAK_EXTERNAL (0x0069)
value IMAGE_SYM_DEBUG ((SHORT)-2)
value IMAGE_SYM_DTYPE_ARRAY (3)
value IMAGE_SYM_DTYPE_FUNCTION (2)
value IMAGE_SYM_DTYPE_NULL (0)
value IMAGE_SYM_DTYPE_POINTER (1)
value IMAGE_SYM_SECTION_MAX (0xFEFF)
value IMAGE_SYM_SECTION_MAX_EX (MAXLONG)
value IMAGE_SYM_TYPE_BYTE (0x000C)
value IMAGE_SYM_TYPE_CHAR (0x0002)
value IMAGE_SYM_TYPE_DOUBLE (0x0007)
value IMAGE_SYM_TYPE_DWORD (0x000F)
value IMAGE_SYM_TYPE_ENUM (0x000A)
value IMAGE_SYM_TYPE_FLOAT (0x0006)
value IMAGE_SYM_TYPE_INT (0x0004)
value IMAGE_SYM_TYPE_LONG (0x0005)
value IMAGE_SYM_TYPE_MOE (0x000B)
value IMAGE_SYM_TYPE_NULL (0x0000)
value IMAGE_SYM_TYPE_PCODE (0x8000)
value IMAGE_SYM_TYPE_SHORT (0x0003)
value IMAGE_SYM_TYPE_STRUCT (0x0008)
value IMAGE_SYM_TYPE_UINT (0x000E)
value IMAGE_SYM_TYPE_UNION (0x0009)
value IMAGE_SYM_TYPE_VOID (0x0001)
value IMAGE_SYM_TYPE_WORD (0x000D)
value IMAGE_SYM_UNDEFINED ((SHORT)0)
value IMAGE_VXD_SIGNATURE (0x454C)
value IMAGE_WEAK_EXTERN_ANTI_DEPENDENCY (4)
value IMAGE_WEAK_EXTERN_SEARCH_ALIAS (3)
value IMAGE_WEAK_EXTERN_SEARCH_LIBRARY (2)
value IMAGE_WEAK_EXTERN_SEARCH_NOLIBRARY (1)
value IMC_CLOSESTATUSWINDOW (0x0021)
value IMC_GETCANDIDATEPOS (0x0007)
value IMC_GETCOMPOSITIONFONT (0x0009)
value IMC_GETCOMPOSITIONWINDOW (0x000B)
value IMC_GETSTATUSWINDOWPOS (0x000F)
value IMC_OPENSTATUSWINDOW (0x0022)
value IMC_SETCANDIDATEPOS (0x0008)
value IMC_SETCOMPOSITIONFONT (0x000A)
value IMC_SETCOMPOSITIONWINDOW (0x000C)
value IMC_SETSTATUSWINDOWPOS (0x0010)
value IMEMENUITEM_STRING_SIZE (80)
value IME_CAND_CODE (0x0002)
value IME_CAND_MEANING (0x0003)
value IME_CAND_RADICAL (0x0004)
value IME_CAND_READ (0x0001)
value IME_CAND_STROKE (0x0005)
value IME_CAND_UNKNOWN (0x0000)
value IME_CHOTKEY_IME_NONIME_TOGGLE (0x10)
value IME_CHOTKEY_SHAPE_TOGGLE (0x11)
value IME_CHOTKEY_SYMBOL_TOGGLE (0x12)
value IME_CMODE_ALPHANUMERIC (0x0000)
value IME_CMODE_CHARCODE (0x0020)
value IME_CMODE_CHINESE (IME_CMODE_NATIVE)
value IME_CMODE_EUDC (0x0200)
value IME_CMODE_FIXED (0x0800)
value IME_CMODE_FULLSHAPE (0x0008)
value IME_CMODE_HANGEUL (IME_CMODE_NATIVE)
value IME_CMODE_HANGUL (IME_CMODE_NATIVE)
value IME_CMODE_HANJACONVERT (0x0040)
value IME_CMODE_JAPANESE (IME_CMODE_NATIVE)
value IME_CMODE_KATAKANA (0x0002)
value IME_CMODE_LANGUAGE (0x0003)
value IME_CMODE_NATIVE (0x0001)
value IME_CMODE_NATIVESYMBOL (0x0080)
value IME_CMODE_NOCONVERSION (0x0100)
value IME_CMODE_RESERVED (0xF0000000)
value IME_CMODE_ROMAN (0x0010)
value IME_CMODE_SOFTKBD (0x0080)
value IME_CMODE_SYMBOL (0x0400)
value IME_CONFIG_GENERAL (1)
value IME_CONFIG_REGISTERWORD (2)
value IME_CONFIG_SELECTDICTIONARY (3)
value IME_ESC_AUTOMATA (0x1009)
value IME_ESC_GETHELPFILENAME (0x100b)
value IME_ESC_GET_EUDC_DICTIONARY (0x1003)
value IME_ESC_HANJA_MODE (0x1008)
value IME_ESC_IME_NAME (0x1006)
value IME_ESC_MAX_KEY (0x1005)
value IME_ESC_PRIVATE_FIRST (0x0800)
value IME_ESC_PRIVATE_HOTKEY (0x100a)
value IME_ESC_PRIVATE_LAST (0x0FFF)
value IME_ESC_QUERY_SUPPORT (0x0003)
value IME_ESC_RESERVED_FIRST (0x0004)
value IME_ESC_RESERVED_LAST (0x07FF)
value IME_ESC_SEQUENCE_TO_INTERNAL (0x1001)
value IME_ESC_SET_EUDC_DICTIONARY (0x1004)
value IME_ESC_SYNC_HOTKEY (0x1007)
value IME_HOTKEY_DSWITCH_FIRST (0x100)
value IME_HOTKEY_DSWITCH_LAST (0x11F)
value IME_HOTKEY_PRIVATE_FIRST (0x200)
value IME_HOTKEY_PRIVATE_LAST (0x21F)
value IME_ITHOTKEY_PREVIOUS_COMPOSITION (0x201)
value IME_ITHOTKEY_RECONVERTSTRING (0x203)
value IME_ITHOTKEY_RESEND_RESULTSTR (0x200)
value IME_ITHOTKEY_UISTYLE_TOGGLE (0x202)
value IME_JHOTKEY_CLOSE_OPEN (0x30)
value IME_KHOTKEY_ENGLISH (0x52)
value IME_KHOTKEY_HANJACONVERT (0x51)
value IME_KHOTKEY_SHAPE_TOGGLE (0x50)
value IME_PROP_AT_CARET (0x00010000)
value IME_PROP_COMPLETE_ON_UNSELECT (0x00100000)
value IME_PROP_SPECIAL_UI (0x00020000)
value IME_PROP_UNICODE (0x00080000)
value IME_REGWORD_STYLE_EUDC (0x00000001)
value IME_REGWORD_STYLE_USER_FIRST (0x80000000)
value IME_REGWORD_STYLE_USER_LAST (0xFFFFFFFF)
value IME_SMODE_AUTOMATIC (0x0004)
value IME_SMODE_CONVERSATION (0x0010)
value IME_SMODE_NONE (0x0000)
value IME_SMODE_PHRASEPREDICT (0x0008)
value IME_SMODE_PLAURALCLAUSE (0x0001)
value IME_SMODE_RESERVED (0x0000F000)
value IME_SMODE_SINGLECONVERT (0x0002)
value IME_THOTKEY_IME_NONIME_TOGGLE (0x70)
value IME_THOTKEY_SHAPE_TOGGLE (0x71)
value IME_THOTKEY_SYMBOL_TOGGLE (0x72)
value IMFS_CHECKED (MFS_CHECKED)
value IMFS_DEFAULT (MFS_DEFAULT)
value IMFS_DISABLED (MFS_DISABLED)
value IMFS_ENABLED (MFS_ENABLED)
value IMFS_GRAYED (MFS_GRAYED)
value IMFS_HILITE (MFS_HILITE)
value IMFS_UNCHECKED (MFS_UNCHECKED)
value IMFS_UNHILITE (MFS_UNHILITE)
value IMFT_RADIOCHECK (0x00001)
value IMFT_SEPARATOR (0x00002)
value IMFT_SUBMENU (0x00004)
value IMM_ERROR_GENERAL ((-2))
value IMM_ERROR_NODATA ((-1))
value IMN_CHANGECANDIDATE (0x0003)
value IMN_CLOSECANDIDATE (0x0004)
value IMN_CLOSESTATUSWINDOW (0x0001)
value IMN_GUIDELINE (0x000D)
value IMN_OPENCANDIDATE (0x0005)
value IMN_OPENSTATUSWINDOW (0x0002)
value IMN_PRIVATE (0x000E)
value IMN_SETCANDIDATEPOS (0x0009)
value IMN_SETCOMPOSITIONFONT (0x000A)
value IMN_SETCOMPOSITIONWINDOW (0x000B)
value IMN_SETCONVERSIONMODE (0x0006)
value IMN_SETOPENSTATUS (0x0008)
value IMN_SETSENTENCEMODE (0x0007)
value IMN_SETSTATUSWINDOWPOS (0x000C)
value IMPLINK_HIGHEXPER (158)
value IMPLINK_IP (155)
value IMPLINK_LOWEXPER (156)
value IMPLTYPEFLAG_FDEFAULT (( 0x1 ))
value IMPLTYPEFLAG_FDEFAULTVTABLE (( 0x8 ))
value IMPLTYPEFLAG_FRESTRICTED (( 0x4 ))
value IMPLTYPEFLAG_FSOURCE (( 0x2 ))
value IMR_CANDIDATEWINDOW (0x0002)
value IMR_COMPOSITIONFONT (0x0003)
value IMR_COMPOSITIONWINDOW (0x0001)
value IMR_CONFIRMRECONVERTSTRING (0x0005)
value IMR_DOCUMENTFEED (0x0007)
value IMR_QUERYCHARPOSITION (0x0006)
value IMR_RECONVERTSTRING (0x0004)
value INADDR_ANY ((ULONG)0x00000000)
value INADDR_LOOPBACK (0x7f000001)
value INADDR_NONE (0xffffffff)
value INCL_WINSOCK_API_PROTOTYPES (1)
value INCL_WINSOCK_API_TYPEDEFS (0)
value INDEXID_CONTAINER (0)
value INDEXID_OBJECT (0)
value INET_E_AUTHENTICATION_REQUIRED (_HRESULT_TYPEDEF_(0x800C0009L))
value INET_E_BLOCKED_ENHANCEDPROTECTEDMODE (_HRESULT_TYPEDEF_(0x800C0506L))
value INET_E_BLOCKED_PLUGGABLE_PROTOCOL (_HRESULT_TYPEDEF_(0x800C0505L))
value INET_E_BLOCKED_REDIRECT_XSECURITYID (_HRESULT_TYPEDEF_(0x800C001BL))
value INET_E_CANNOT_CONNECT (_HRESULT_TYPEDEF_(0x800C0004L))
value INET_E_CANNOT_INSTANTIATE_OBJECT (_HRESULT_TYPEDEF_(0x800C0010L))
value INET_E_CANNOT_LOAD_DATA (_HRESULT_TYPEDEF_(0x800C000FL))
value INET_E_CANNOT_LOCK_REQUEST (_HRESULT_TYPEDEF_(0x800C0016L))
value INET_E_CANNOT_REPLACE_SFP_FILE (_HRESULT_TYPEDEF_(0x800C0300L))
value INET_E_CODE_DOWNLOAD_DECLINED (_HRESULT_TYPEDEF_(0x800C0100L))
value INET_E_CODE_INSTALL_BLOCKED_ARM (_HRESULT_TYPEDEF_(0x800C0504L))
value INET_E_CODE_INSTALL_BLOCKED_BITNESS (_HRESULT_TYPEDEF_(0x800C0507L))
value INET_E_CODE_INSTALL_BLOCKED_BY_HASH_POLICY (_HRESULT_TYPEDEF_(0x800C0500L))
value INET_E_CODE_INSTALL_BLOCKED_IMMERSIVE (_HRESULT_TYPEDEF_(0x800C0502L))
value INET_E_CODE_INSTALL_SUPPRESSED (_HRESULT_TYPEDEF_(0x800C0400L))
value INET_E_CONNECTION_TIMEOUT (_HRESULT_TYPEDEF_(0x800C000BL))
value INET_E_DATA_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x800C0007L))
value INET_E_DEFAULT_ACTION (INET_E_USE_DEFAULT_PROTOCOLHANDLER)
value INET_E_DOMINJECTIONVALIDATION (_HRESULT_TYPEDEF_(0x800C001CL))
value INET_E_DOWNLOAD_BLOCKED_BY_CSP (_HRESULT_TYPEDEF_(0x800C0508L))
value INET_E_DOWNLOAD_BLOCKED_BY_INPRIVATE (_HRESULT_TYPEDEF_(0x800C0501L))
value INET_E_DOWNLOAD_FAILURE (_HRESULT_TYPEDEF_(0x800C0008L))
value INET_E_ERROR_FIRST (_HRESULT_TYPEDEF_(0x800C0002L))
value INET_E_ERROR_LAST (INET_E_DOWNLOAD_BLOCKED_BY_CSP)
value INET_E_FORBIDFRAMING (_HRESULT_TYPEDEF_(0x800C0503L))
value INET_E_HSTS_CERTIFICATE_ERROR (_HRESULT_TYPEDEF_(0x800C001EL))
value INET_E_INVALID_CERTIFICATE (_HRESULT_TYPEDEF_(0x800C0019L))
value INET_E_INVALID_REQUEST (_HRESULT_TYPEDEF_(0x800C000CL))
value INET_E_INVALID_URL (_HRESULT_TYPEDEF_(0x800C0002L))
value INET_E_NO_SESSION (_HRESULT_TYPEDEF_(0x800C0003L))
value INET_E_NO_VALID_MEDIA (_HRESULT_TYPEDEF_(0x800C000AL))
value INET_E_OBJECT_NOT_FOUND (_HRESULT_TYPEDEF_(0x800C0006L))
value INET_E_QUERYOPTION_UNKNOWN (_HRESULT_TYPEDEF_(0x800C0013L))
value INET_E_REDIRECTING (_HRESULT_TYPEDEF_(0x800C0014L))
value INET_E_REDIRECT_FAILED (_HRESULT_TYPEDEF_(0x800C0014L))
value INET_E_REDIRECT_TO_DIR (_HRESULT_TYPEDEF_(0x800C0015L))
value INET_E_RESOURCE_NOT_FOUND (_HRESULT_TYPEDEF_(0x800C0005L))
value INET_E_RESULT_DISPATCHED (_HRESULT_TYPEDEF_(0x800C0200L))
value INET_E_SECURITY_PROBLEM (_HRESULT_TYPEDEF_(0x800C000EL))
value INET_E_TERMINATED_BIND (_HRESULT_TYPEDEF_(0x800C0018L))
value INET_E_UNKNOWN_PROTOCOL (_HRESULT_TYPEDEF_(0x800C000DL))
value INET_E_USE_DEFAULT_PROTOCOLHANDLER (_HRESULT_TYPEDEF_(0x800C0011L))
value INET_E_USE_DEFAULT_SETTING (_HRESULT_TYPEDEF_(0x800C0012L))
value INET_E_USE_EXTEND_BINDING (_HRESULT_TYPEDEF_(0x800C0017L))
value INET_E_VTAB_SWITCH_FORCE_ENGINE (_HRESULT_TYPEDEF_(0x800C001DL))
value INFINITE (0xFFFFFFFF)
value INHERITED_ACE ((0x10))
value INHERIT_CALLER_PRIORITY (0x00020000)
value INHERIT_ONLY_ACE ((0x8))
value INHERIT_PARENT_AFFINITY (0x00010000)
value INITIAL_FPCSR (0x027f)
value INITIAL_MXCSR (0x1f80)
value INIT_ONCE_ASYNC (RTL_RUN_ONCE_ASYNC)
value INIT_ONCE_CHECK_ONLY (RTL_RUN_ONCE_CHECK_ONLY)
value INIT_ONCE_CTX_RESERVED_BITS (RTL_RUN_ONCE_CTX_RESERVED_BITS)
value INIT_ONCE_INIT_FAILED (RTL_RUN_ONCE_INIT_FAILED)
value INIT_ONCE_STATIC_INIT (RTL_RUN_ONCE_INIT)
value INPLACE_E_FIRST (0x800401A0L)
value INPLACE_E_LAST (0x800401AFL)
value INPLACE_E_NOTOOLSPACE (_HRESULT_TYPEDEF_(0x800401A1L))
value INPLACE_E_NOTUNDOABLE (_HRESULT_TYPEDEF_(0x800401A0L))
value INPLACE_S_FIRST (0x000401A0L)
value INPLACE_S_LAST (0x000401AFL)
value INPLACE_S_TRUNCATED (_HRESULT_TYPEDEF_(0x000401A0L))
value INPUTLANGCHANGE_BACKWARD (0x0004)
value INPUTLANGCHANGE_FORWARD (0x0002)
value INPUTLANGCHANGE_SYSCHARSET (0x0001)
value INPUT_E_DEVICE_INFO (_HRESULT_TYPEDEF_(0x80400006L))
value INPUT_E_DEVICE_PROPERTY (_HRESULT_TYPEDEF_(0x80400008L))
value INPUT_E_FRAME (_HRESULT_TYPEDEF_(0x80400004L))
value INPUT_E_HISTORY (_HRESULT_TYPEDEF_(0x80400005L))
value INPUT_E_MULTIMODAL (_HRESULT_TYPEDEF_(0x80400002L))
value INPUT_E_OUT_OF_ORDER (_HRESULT_TYPEDEF_(0x80400000L))
value INPUT_E_PACKET (_HRESULT_TYPEDEF_(0x80400003L))
value INPUT_E_REENTRANCY (_HRESULT_TYPEDEF_(0x80400001L))
value INPUT_E_TRANSFORM (_HRESULT_TYPEDEF_(0x80400007L))
value INPUT_HARDWARE (2)
value INPUT_KEYBOARD (1)
value INPUT_MOUSE (0)
value INTERNATIONAL_USAGE (0x00000001)
value INT_MAX (2147483647)
value INT_MIN ((-2147483647 - 1))
value INVALID_ATOM (((ATOM)0))
value INVALID_FILE_ATTRIBUTES (((DWORD)-1))
value INVALID_FILE_SIZE (((DWORD)0xFFFFFFFF))
value INVALID_HANDLE_VALUE (((HANDLE)(LONG_PTR)-1))
value INVALID_SET_FILE_POINTER (((DWORD)-1))
value IN_CLASSA_HOST (0x00ffffff)
value IN_CLASSA_MAX (128)
value IN_CLASSA_NET (0xff000000)
value IN_CLASSA_NSHIFT (24)
value IN_CLASSB_HOST (0x0000ffff)
value IN_CLASSB_MAX (65536)
value IN_CLASSB_NET (0xffff0000)
value IN_CLASSB_NSHIFT (16)
value IN_CLASSC_HOST (0x000000ff)
value IN_CLASSC_NET (0xffffff00)
value IN_CLASSC_NSHIFT (8)
value IN_CLASSD_HOST (0x0fffffff)
value IN_CLASSD_NET (0xf0000000)
value IN_CLASSD_NSHIFT (28)
value IOCPARM_MASK (0x7f)
value IOCTL_CHANGER_BASE (FILE_DEVICE_CHANGER)
value IOCTL_DISK_BASE (FILE_DEVICE_DISK)
value IOCTL_SCMBUS_BASE (FILE_DEVICE_PERSISTENT_MEMORY)
value IOCTL_SCMBUS_DEVICE_FUNCTION_BASE (0x0)
value IOCTL_SCM_LOGICAL_DEVICE_FUNCTION_BASE (0x300)
value IOCTL_SCM_PHYSICAL_DEVICE_FUNCTION_BASE (0x600)
value IOCTL_SMARTCARD_CONFISCATE (SCARD_CTL_CODE( 4))
value IOCTL_SMARTCARD_EJECT (SCARD_CTL_CODE( 6))
value IOCTL_SMARTCARD_GET_ATTRIBUTE (SCARD_CTL_CODE( 2))
value IOCTL_SMARTCARD_GET_FEATURE_REQUEST (SCARD_CTL_CODE(3400))
value IOCTL_SMARTCARD_GET_LAST_ERROR (SCARD_CTL_CODE(15))
value IOCTL_SMARTCARD_GET_PERF_CNTR (SCARD_CTL_CODE(16))
value IOCTL_SMARTCARD_GET_STATE (SCARD_CTL_CODE(14))
value IOCTL_SMARTCARD_IS_ABSENT (SCARD_CTL_CODE(11))
value IOCTL_SMARTCARD_IS_PRESENT (SCARD_CTL_CODE(10))
value IOCTL_SMARTCARD_POWER (SCARD_CTL_CODE( 1))
value IOCTL_SMARTCARD_SET_ATTRIBUTE (SCARD_CTL_CODE( 3))
value IOCTL_SMARTCARD_SET_PROTOCOL (SCARD_CTL_CODE(12))
value IOCTL_SMARTCARD_SWALLOW (SCARD_CTL_CODE( 7))
value IOCTL_SMARTCARD_TRANSMIT (SCARD_CTL_CODE( 5))
value IOCTL_STORAGE_BASE (FILE_DEVICE_MASS_STORAGE)
value IOCTL_STORAGE_BC_VERSION (1)
value IOCTL_VOLUME_BASE (0x00000056)
value IOC_IN (0x80000000)
value IOC_INOUT ((IOC_IN|IOC_OUT))
value IOC_OUT (0x40000000)
value IOC_PROTOCOL (0x10000000)
value IOC_UNIX (0x00000000)
value IOC_VENDOR (0x18000000)
value IOC_VOID (0x20000000)
value IOC_WSK ((IOC_WS2|0x07000000))
value IORING_E_COMPLETION_QUEUE_TOO_BIG (_HRESULT_TYPEDEF_(0x80460005L))
value IORING_E_COMPLETION_QUEUE_TOO_FULL (_HRESULT_TYPEDEF_(0x80460008L))
value IORING_E_CORRUPT (_HRESULT_TYPEDEF_(0x80460007L))
value IORING_E_REQUIRED_FLAG_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80460001L))
value IORING_E_SUBMISSION_QUEUE_FULL (_HRESULT_TYPEDEF_(0x80460002L))
value IORING_E_SUBMISSION_QUEUE_TOO_BIG (_HRESULT_TYPEDEF_(0x80460004L))
value IORING_E_SUBMIT_IN_PROGRESS (_HRESULT_TYPEDEF_(0x80460006L))
value IORING_E_VERSION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80460003L))
value IO_COMPLETION_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED|SYNCHRONIZE|0x3))
value IO_COMPLETION_MODIFY_STATE (0x0002)
value IO_QOS_MAX_RESERVATION (1000000000ULL)
value IO_REPARSE_TAG_AF_UNIX ((0x80000023L))
value IO_REPARSE_TAG_APPEXECLINK ((0x8000001BL))
value IO_REPARSE_TAG_CLOUD ((0x9000001AL))
value IO_REPARSE_TAG_CLOUD_A ((0x9000A01AL))
value IO_REPARSE_TAG_CLOUD_B ((0x9000B01AL))
value IO_REPARSE_TAG_CLOUD_C ((0x9000C01AL))
value IO_REPARSE_TAG_CLOUD_D ((0x9000D01AL))
value IO_REPARSE_TAG_CLOUD_E ((0x9000E01AL))
value IO_REPARSE_TAG_CLOUD_F ((0x9000F01AL))
value IO_REPARSE_TAG_CLOUD_MASK ((0x0000F000L))
value IO_REPARSE_TAG_CSV ((0x80000009L))
value IO_REPARSE_TAG_DATALESS_CIM ((0xA0000028L))
value IO_REPARSE_TAG_DEDUP ((0x80000013L))
value IO_REPARSE_TAG_DFS ((0x8000000AL))
value IO_REPARSE_TAG_DFSR ((0x80000012L))
value IO_REPARSE_TAG_FILE_PLACEHOLDER ((0x80000015L))
value IO_REPARSE_TAG_GLOBAL_REPARSE ((0xA0000019L))
value IO_REPARSE_TAG_HSM ((0xC0000004L))
value IO_REPARSE_TAG_MOUNT_POINT ((0xA0000003L))
value IO_REPARSE_TAG_NFS ((0x80000014L))
value IO_REPARSE_TAG_ONEDRIVE ((0x80000021L))
value IO_REPARSE_TAG_PROJFS ((0x9000001CL))
value IO_REPARSE_TAG_PROJFS_TOMBSTONE ((0xA0000022L))
value IO_REPARSE_TAG_RESERVED_ONE ((1))
value IO_REPARSE_TAG_RESERVED_RANGE (IO_REPARSE_TAG_RESERVED_TWO)
value IO_REPARSE_TAG_RESERVED_TWO ((2))
value IO_REPARSE_TAG_RESERVED_ZERO ((0))
value IO_REPARSE_TAG_SIS ((0x80000007L))
value IO_REPARSE_TAG_STORAGE_SYNC ((0x8000001EL))
value IO_REPARSE_TAG_SYMLINK ((0xA000000CL))
value IO_REPARSE_TAG_UNHANDLED ((0x80000020L))
value IO_REPARSE_TAG_WCI ((0x80000018L))
value IO_REPARSE_TAG_WCI_LINK ((0xA0000027L))
value IO_REPARSE_TAG_WCI_TOMBSTONE ((0xA000001FL))
value IO_REPARSE_TAG_WIM ((0x80000008L))
value IO_REPARSE_TAG_WOF ((0x80000017L))
value IPDFP_COPY_ALL_FILES (0x00000001)
value IPPORT_BIFFUDP (512)
value IPPORT_CHARGEN (19)
value IPPORT_CMDSERVER (514)
value IPPORT_DAYTIME (13)
value IPPORT_DISCARD (9)
value IPPORT_DYNAMIC_MAX (0xffff)
value IPPORT_DYNAMIC_MIN (0xc000)
value IPPORT_ECHO (7)
value IPPORT_EFSSERVER (520)
value IPPORT_EPMAP (135)
value IPPORT_EXECSERVER (512)
value IPPORT_FINGER (79)
value IPPORT_FTP (21)
value IPPORT_FTP_DATA (20)
value IPPORT_HTTPS (443)
value IPPORT_IMAP (143)
value IPPORT_LDAP (389)
value IPPORT_LOGINSERVER (513)
value IPPORT_MICROSOFT_DS (445)
value IPPORT_MSP (18)
value IPPORT_MTP (57)
value IPPORT_NAMESERVER (42)
value IPPORT_NETBIOS_DGM (138)
value IPPORT_NETBIOS_NS (137)
value IPPORT_NETBIOS_SSN (139)
value IPPORT_NETSTAT (15)
value IPPORT_NTP (123)
value IPPORT_QOTD (17)
value IPPORT_REGISTERED_MAX (0xbfff)
value IPPORT_REGISTERED_MIN (IPPORT_RESERVED)
value IPPORT_RESERVED (1024)
value IPPORT_RJE (77)
value IPPORT_ROUTESERVER (520)
value IPPORT_SMTP (25)
value IPPORT_SNMP (161)
value IPPORT_SNMP_TRAP (162)
value IPPORT_SUPDUP (95)
value IPPORT_SYSTAT (11)
value IPPORT_TCPMUX (1)
value IPPORT_TELNET (23)
value IPPORT_TFTP (69)
value IPPORT_TIMESERVER (37)
value IPPORT_TTYLINK (87)
value IPPORT_WHOIS (43)
value IPPORT_WHOSERVER (513)
value IPPROTO_IP (0)
value ISC_SHOWUIALL (0xC000000F)
value ISC_SHOWUIALLCANDIDATEWINDOW (0x0000000F)
value ISC_SHOWUICANDIDATEWINDOW (0x00000001)
value ISC_SHOWUICOMPOSITIONWINDOW (0x80000000)
value ISC_SHOWUIGUIDELINE (0x40000000)
value ISMEX_CALLBACK (0x00000004)
value ISMEX_NOSEND (0x00000000)
value ISMEX_NOTIFY (0x00000002)
value ISMEX_REPLIED (0x00000008)
value ISMEX_SEND (0x00000001)
value ISOLATIONAWARE_MANIFEST_RESOURCE_ID (MAKEINTRESOURCE(2))
value ISOLATIONAWARE_NOSTATICIMPORT_MANIFEST_RESOURCE_ID (MAKEINTRESOURCE(3))
value ISOLATIONPOLICY_BROWSER_MANIFEST_RESOURCE_ID (MAKEINTRESOURCE(5))
value ISOLATIONPOLICY_MANIFEST_RESOURCE_ID (MAKEINTRESOURCE(4))
value IS_TEXT_UNICODE_CONTROLS (0x0004)
value IS_TEXT_UNICODE_DBCS_LEADBYTE (0x0400)
value IS_TEXT_UNICODE_ILLEGAL_CHARS (0x0100)
value IS_TEXT_UNICODE_NOT_ASCII_MASK (0xF000)
value IS_TEXT_UNICODE_NOT_UNICODE_MASK (0x0F00)
value IS_TEXT_UNICODE_NULL_BYTES (0x1000)
value IS_TEXT_UNICODE_ODD_LENGTH (0x0200)
value IS_TEXT_UNICODE_REVERSE_CONTROLS (0x0040)
value IS_TEXT_UNICODE_REVERSE_MASK (0x00F0)
value IS_TEXT_UNICODE_REVERSE_SIGNATURE (0x0080)
value IS_TEXT_UNICODE_REVERSE_STATISTICS (0x0020)
value IS_TEXT_UNICODE_SIGNATURE (0x0008)
value IS_TEXT_UNICODE_STATISTICS (0x0002)
value IS_TEXT_UNICODE_UNICODE_MASK (0x000F)
value ITALIC_FONTTYPE (0x0200)
value I_RRPCUNINITIALIZENDROLE_EXPORT_NAME (((LPCSTR)(ULONG_PTR)1000))
value JL_BOTH (0x04)
value JL_RECEIVER_ONLY (0x02)
value JL_SENDER_ONLY (0x01)
value JOB_ACCESS_ADMINISTER (0x00000010)
value JOB_ACCESS_READ (0x00000020)
value JOB_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | JOB_ACCESS_ADMINISTER | JOB_ACCESS_READ))
value JOB_CONTROL_CANCEL (3)
value JOB_CONTROL_DELETE (5)
value JOB_CONTROL_LAST_PAGE_EJECTED (7)
value JOB_CONTROL_PAUSE (1)
value JOB_CONTROL_RELEASE (9)
value JOB_CONTROL_RESTART (4)
value JOB_CONTROL_RESUME (2)
value JOB_CONTROL_RETAIN (8)
value JOB_CONTROL_SEND_TOAST (10)
value JOB_CONTROL_SENT_TO_PRINTER (6)
value JOB_EXECUTE ((STANDARD_RIGHTS_EXECUTE | JOB_ACCESS_ADMINISTER))
value JOB_NOTIFY_FIELD_BYTES_PRINTED (0x17)
value JOB_NOTIFY_FIELD_DATATYPE (0x05)
value JOB_NOTIFY_FIELD_DEVMODE (0x09)
value JOB_NOTIFY_FIELD_DOCUMENT (0x0D)
value JOB_NOTIFY_FIELD_DRIVER_NAME (0x08)
value JOB_NOTIFY_FIELD_MACHINE_NAME (0x01)
value JOB_NOTIFY_FIELD_NOTIFY_NAME (0x04)
value JOB_NOTIFY_FIELD_PAGES_PRINTED (0x15)
value JOB_NOTIFY_FIELD_PARAMETERS (0x07)
value JOB_NOTIFY_FIELD_PORT_NAME (0x02)
value JOB_NOTIFY_FIELD_POSITION (0x0F)
value JOB_NOTIFY_FIELD_PRINTER_NAME (0x00)
value JOB_NOTIFY_FIELD_PRINT_PROCESSOR (0x06)
value JOB_NOTIFY_FIELD_PRIORITY (0x0E)
value JOB_NOTIFY_FIELD_REMOTE_JOB_ID (0x18)
value JOB_NOTIFY_FIELD_SECURITY_DESCRIPTOR (0x0C)
value JOB_NOTIFY_FIELD_START_TIME (0x11)
value JOB_NOTIFY_FIELD_STATUS (0x0A)
value JOB_NOTIFY_FIELD_STATUS_STRING (0x0B)
value JOB_NOTIFY_FIELD_SUBMITTED (0x10)
value JOB_NOTIFY_FIELD_TIME (0x13)
value JOB_NOTIFY_FIELD_TOTAL_BYTES (0x16)
value JOB_NOTIFY_FIELD_TOTAL_PAGES (0x14)
value JOB_NOTIFY_FIELD_UNTIL_TIME (0x12)
value JOB_NOTIFY_FIELD_USER_NAME (0x03)
value JOB_NOTIFY_TYPE (0x01)
value JOB_OBJECT_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | SYNCHRONIZE | 0x3F ))
value JOB_OBJECT_ASSIGN_PROCESS ((0x0001))
value JOB_OBJECT_BASIC_LIMIT_VALID_FLAGS (0x000000ff)
value JOB_OBJECT_CPU_RATE_CONTROL_ENABLE (0x1)
value JOB_OBJECT_CPU_RATE_CONTROL_HARD_CAP (0x4)
value JOB_OBJECT_CPU_RATE_CONTROL_MIN_MAX_RATE (0x10)
value JOB_OBJECT_CPU_RATE_CONTROL_NOTIFY (0x8)
value JOB_OBJECT_CPU_RATE_CONTROL_VALID_FLAGS (0x1f)
value JOB_OBJECT_CPU_RATE_CONTROL_WEIGHT_BASED (0x2)
value JOB_OBJECT_EXTENDED_LIMIT_VALID_FLAGS (0x00007fff)
value JOB_OBJECT_IMPERSONATE ((0x0020))
value JOB_OBJECT_LIMIT_ACTIVE_PROCESS (0x00000008)
value JOB_OBJECT_LIMIT_AFFINITY (0x00000010)
value JOB_OBJECT_LIMIT_BREAKAWAY_OK (0x00000800)
value JOB_OBJECT_LIMIT_CPU_RATE_CONTROL (JOB_OBJECT_LIMIT_RATE_CONTROL)
value JOB_OBJECT_LIMIT_DIE_ON_UNHANDLED_EXCEPTION (0x00000400)
value JOB_OBJECT_LIMIT_IO_RATE_CONTROL (0x00080000)
value JOB_OBJECT_LIMIT_JOB_MEMORY (0x00000200)
value JOB_OBJECT_LIMIT_JOB_MEMORY_HIGH (JOB_OBJECT_LIMIT_JOB_MEMORY)
value JOB_OBJECT_LIMIT_JOB_MEMORY_LOW (0x00008000)
value JOB_OBJECT_LIMIT_JOB_READ_BYTES (0x00010000)
value JOB_OBJECT_LIMIT_JOB_TIME (0x00000004)
value JOB_OBJECT_LIMIT_JOB_WRITE_BYTES (0x00020000)
value JOB_OBJECT_LIMIT_KILL_ON_JOB_CLOSE (0x00002000)
value JOB_OBJECT_LIMIT_NET_RATE_CONTROL (0x00100000)
value JOB_OBJECT_LIMIT_PRESERVE_JOB_TIME (0x00000040)
value JOB_OBJECT_LIMIT_PRIORITY_CLASS (0x00000020)
value JOB_OBJECT_LIMIT_PROCESS_MEMORY (0x00000100)
value JOB_OBJECT_LIMIT_PROCESS_TIME (0x00000002)
value JOB_OBJECT_LIMIT_RATE_CONTROL (0x00040000)
value JOB_OBJECT_LIMIT_SCHEDULING_CLASS (0x00000080)
value JOB_OBJECT_LIMIT_SILENT_BREAKAWAY_OK (0x00001000)
value JOB_OBJECT_LIMIT_SUBSET_AFFINITY (0x00004000)
value JOB_OBJECT_LIMIT_VALID_FLAGS (0x0007ffff)
value JOB_OBJECT_LIMIT_WORKINGSET (0x00000001)
value JOB_OBJECT_MSG_ABNORMAL_EXIT_PROCESS (8)
value JOB_OBJECT_MSG_ACTIVE_PROCESS_LIMIT (3)
value JOB_OBJECT_MSG_ACTIVE_PROCESS_ZERO (4)
value JOB_OBJECT_MSG_END_OF_JOB_TIME (1)
value JOB_OBJECT_MSG_END_OF_PROCESS_TIME (2)
value JOB_OBJECT_MSG_EXIT_PROCESS (7)
value JOB_OBJECT_MSG_JOB_CYCLE_TIME_LIMIT (12)
value JOB_OBJECT_MSG_JOB_MEMORY_LIMIT (10)
value JOB_OBJECT_MSG_MAXIMUM (13)
value JOB_OBJECT_MSG_MINIMUM (1)
value JOB_OBJECT_MSG_NEW_PROCESS (6)
value JOB_OBJECT_MSG_NOTIFICATION_LIMIT (11)
value JOB_OBJECT_MSG_PROCESS_MEMORY_LIMIT (9)
value JOB_OBJECT_MSG_SILO_TERMINATED (13)
value JOB_OBJECT_NET_RATE_CONTROL_MAX_DSCP_TAG (64)
value JOB_OBJECT_NOTIFICATION_LIMIT_VALID_FLAGS ((JOB_OBJECT_LIMIT_JOB_READ_BYTES | JOB_OBJECT_LIMIT_JOB_WRITE_BYTES | JOB_OBJECT_LIMIT_JOB_TIME | JOB_OBJECT_LIMIT_JOB_MEMORY_LOW | JOB_OBJECT_LIMIT_JOB_MEMORY_HIGH | JOB_OBJECT_LIMIT_CPU_RATE_CONTROL | JOB_OBJECT_LIMIT_IO_RATE_CONTROL | JOB_OBJECT_LIMIT_NET_RATE_CONTROL))
value JOB_OBJECT_POST_AT_END_OF_JOB (1)
value JOB_OBJECT_QUERY ((0x0004))
value JOB_OBJECT_SECURITY_FILTER_TOKENS (0x00000008)
value JOB_OBJECT_SECURITY_NO_ADMIN (0x00000001)
value JOB_OBJECT_SECURITY_ONLY_TOKEN (0x00000004)
value JOB_OBJECT_SECURITY_RESTRICTED_TOKEN (0x00000002)
value JOB_OBJECT_SECURITY_VALID_FLAGS (0x0000000f)
value JOB_OBJECT_SET_ATTRIBUTES ((0x0002))
value JOB_OBJECT_SET_SECURITY_ATTRIBUTES ((0x0010))
value JOB_OBJECT_TERMINATE ((0x0008))
value JOB_OBJECT_TERMINATE_AT_END_OF_JOB (0)
value JOB_OBJECT_UILIMIT_ALL (0x000001FF)
value JOB_OBJECT_UILIMIT_DESKTOP (0x00000040)
value JOB_OBJECT_UILIMIT_DISPLAYSETTINGS (0x00000010)
value JOB_OBJECT_UILIMIT_EXITWINDOWS (0x00000080)
value JOB_OBJECT_UILIMIT_GLOBALATOMS (0x00000020)
value JOB_OBJECT_UILIMIT_HANDLES (0x00000001)
value JOB_OBJECT_UILIMIT_IME (0x00000100)
value JOB_OBJECT_UILIMIT_NONE (0x00000000)
value JOB_OBJECT_UILIMIT_READCLIPBOARD (0x00000002)
value JOB_OBJECT_UILIMIT_SYSTEMPARAMETERS (0x00000008)
value JOB_OBJECT_UILIMIT_WRITECLIPBOARD (0x00000004)
value JOB_OBJECT_UI_VALID_FLAGS (0x000001FF)
value JOB_POSITION_UNSPECIFIED (0)
value JOB_READ ((STANDARD_RIGHTS_READ | JOB_ACCESS_READ))
value JOB_STATUS_BLOCKED_DEVQ (0x00000200)
value JOB_STATUS_COMPLETE (0x00001000)
value JOB_STATUS_DELETED (0x00000100)
value JOB_STATUS_DELETING (0x00000004)
value JOB_STATUS_ERROR (0x00000002)
value JOB_STATUS_OFFLINE (0x00000020)
value JOB_STATUS_PAPEROUT (0x00000040)
value JOB_STATUS_PAUSED (0x00000001)
value JOB_STATUS_PRINTED (0x00000080)
value JOB_STATUS_PRINTING (0x00000010)
value JOB_STATUS_RENDERING_LOCALLY (0x00004000)
value JOB_STATUS_RESTART (0x00000800)
value JOB_STATUS_RETAINED (0x00002000)
value JOB_STATUS_SPOOLING (0x00000008)
value JOB_STATUS_USER_INTERVENTION (0x00000400)
value JOB_WRITE ((STANDARD_RIGHTS_WRITE | JOB_ACCESS_ADMINISTER))
value JOHAB_CHARSET (130)
value JOYCAPS_HASPOV (0x0010)
value JOYCAPS_HASR (0x0002)
value JOYCAPS_HASU (0x0004)
value JOYCAPS_HASV (0x0008)
value JOYCAPS_HASZ (0x0001)
value JOYCAPS_POVCTS (0x0040)
value JOYERR_BASE (160)
value JOYERR_NOCANDO ((JOYERR_BASE+6))
value JOYERR_NOERROR ((0))
value JOYERR_PARMS ((JOYERR_BASE+5))
value JOYERR_UNPLUGGED ((JOYERR_BASE+7))
value JOY_POVBACKWARD (18000)
value JOY_POVCENTERED ((WORD) -1)
value JOY_POVFORWARD (0)
value JOY_POVLEFT (27000)
value JOY_POVRIGHT (9000)
value JOY_RETURNALL ((JOY_RETURNX | JOY_RETURNY | JOY_RETURNZ | JOY_RETURNR | JOY_RETURNU | JOY_RETURNV | JOY_RETURNPOV | JOY_RETURNBUTTONS))
value JSCRIPT_E_CANTEXECUTE (_HRESULT_TYPEDEF_(0x89020001L))
value KDF_ALGORITHMID (0x8)
value KDF_CONTEXT (0xE)
value KDF_GENERIC_PARAMETER (0x11)
value KDF_HASH_ALGORITHM (0x0)
value KDF_HKDF_INFO (0x14)
value KDF_HKDF_SALT (0x13)
value KDF_HMAC_KEY (0x3)
value KDF_ITERATION_COUNT (0x10)
value KDF_KEYBITLENGTH (0x12)
value KDF_LABEL (0xD)
value KDF_PARTYUINFO (0x9)
value KDF_PARTYVINFO (0xA)
value KDF_SALT (0xF)
value KDF_SECRET_APPEND (0x2)
value KDF_SECRET_HANDLE (0x6)
value KDF_SECRET_PREPEND (0x1)
value KDF_SUPPPRIVINFO (0xC)
value KDF_SUPPPUBINFO (0xB)
value KDF_TLS_PRF_LABEL (0x4)
value KDF_TLS_PRF_PROTOCOL (0x7)
value KDF_TLS_PRF_SEED (0x5)
value KDF_USE_SECRET_AS_HMAC_KEY_FLAG (0x1)
value KEYBOARD_OVERRUN_MAKE_CODE (0xFF)
value KEYEVENTF_EXTENDEDKEY (0x0001)
value KEYEVENTF_KEYUP (0x0002)
value KEYEVENTF_SCANCODE (0x0008)
value KEYEVENTF_UNICODE (0x0004)
value KEYSTATEBLOB (0xC)
value KEY_CREATE_LINK ((0x0020))
value KEY_CREATE_SUB_KEY ((0x0004))
value KEY_ENUMERATE_SUB_KEYS ((0x0008))
value KEY_EVENT (0x0001)
value KEY_LENGTH_MASK (0xFFFF0000)
value KEY_NOTIFY ((0x0010))
value KEY_QUERY_VALUE ((0x0001))
value KEY_SET_VALUE ((0x0002))
value KF_ALTDOWN (0x2000)
value KF_DLGMODE (0x0800)
value KF_EXTENDED (0x0100)
value KF_MENUMODE (0x1000)
value KF_REPEAT (0x4000)
value KF_UP (0x8000)
value KLF_ACTIVATE (0x00000001)
value KLF_NOTELLSHELL (0x00000080)
value KLF_REORDER (0x00000008)
value KLF_REPLACELANG (0x00000010)
value KLF_RESET (0x40000000)
value KLF_SETFORPROCESS (0x00000100)
value KLF_SHIFTLOCK (0x00010000)
value KLF_SUBSTITUTE_OK (0x00000002)
value KL_NAMELENGTH (9)
value KP_ADMIN_PIN (31)
value KP_ALGID (7)
value KP_BLOCKLEN (8)
value KP_CERTIFICATE (26)
value KP_CLEAR_KEY (27)
value KP_CLIENT_RANDOM (21)
value KP_CMS_DH_KEY_INFO (38)
value KP_CMS_KEY_INFO (37)
value KP_EFFECTIVE_KEYLEN (19)
value KP_G (12)
value KP_GET_USE_COUNT (42)
value KP_HIGHEST_VERSION (41)
value KP_INFO (18)
value KP_IV (1)
value KP_KEYEXCHANGE_PIN (32)
value KP_KEYLEN (9)
value KP_KEYVAL (30)
value KP_MODE (4)
value KP_MODE_BITS (5)
value KP_OAEP_PARAMS (36)
value KP_P (11)
value KP_PADDING (3)
value KP_PERMISSIONS (6)
value KP_PIN_ID (43)
value KP_PIN_INFO (44)
value KP_PRECOMP_SHA (25)
value KP_PREHASH (34)
value KP_PUB_EX_LEN (28)
value KP_PUB_EX_VAL (29)
value KP_PUB_PARAMS (39)
value KP_Q (13)
value KP_RA (16)
value KP_RB (17)
value KP_ROUNDS (35)
value KP_RP (23)
value KP_SALT (2)
value KP_SALT_EX (10)
value KP_SCHANNEL_ALG (20)
value KP_SERVER_RANDOM (22)
value KP_SIGNATURE_PIN (33)
value KP_VERIFY_PARAMS (40)
value KP_X (14)
value KP_Y (15)
value KTM_MARSHAL_BLOB_VERSION_MAJOR (1)
value KTM_MARSHAL_BLOB_VERSION_MINOR (1)
value LABEL_SECURITY_INFORMATION ((0x00000010L))
value LANGGROUPLOCALE_ENUMPROC (LANGGROUPLOCALE_ENUMPROCA)
value LANGUAGEGROUP_ENUMPROC (LANGUAGEGROUP_ENUMPROCA)
value LANG_AFRIKAANS (0x36)
value LANG_ALBANIAN (0x1c)
value LANG_ALSATIAN (0x84)
value LANG_AMHARIC (0x5e)
value LANG_ARABIC (0x01)
value LANG_ARMENIAN (0x2b)
value LANG_ASSAMESE (0x4d)
value LANG_AZERBAIJANI (0x2c)
value LANG_AZERI (0x2c)
value LANG_BANGLA (0x45)
value LANG_BASHKIR (0x6d)
value LANG_BASQUE (0x2d)
value LANG_BELARUSIAN (0x23)
value LANG_BENGALI (0x45)
value LANG_BOSNIAN (0x1a)
value LANG_BOSNIAN_NEUTRAL (0x781a)
value LANG_BRETON (0x7e)
value LANG_BULGARIAN (0x02)
value LANG_CATALAN (0x03)
value LANG_CENTRAL_KURDISH (0x92)
value LANG_CHEROKEE (0x5c)
value LANG_CHINESE (0x04)
value LANG_CHINESE_SIMPLIFIED (0x04)
value LANG_CHINESE_TRADITIONAL (0x7c04)
value LANG_CORSICAN (0x83)
value LANG_CROATIAN (0x1a)
value LANG_CZECH (0x05)
value LANG_DANISH (0x06)
value LANG_DARI (0x8c)
value LANG_DIVEHI (0x65)
value LANG_DUTCH (0x13)
value LANG_ENGLISH (0x09)
value LANG_ESTONIAN (0x25)
value LANG_FAEROESE (0x38)
value LANG_FARSI (0x29)
value LANG_FILIPINO (0x64)
value LANG_FINNISH (0x0b)
value LANG_FRENCH (0x0c)
value LANG_FRISIAN (0x62)
value LANG_FULAH (0x67)
value LANG_GALICIAN (0x56)
value LANG_GEORGIAN (0x37)
value LANG_GERMAN (0x07)
value LANG_GREEK (0x08)
value LANG_GREENLANDIC (0x6f)
value LANG_GUJARATI (0x47)
value LANG_HAUSA (0x68)
value LANG_HAWAIIAN (0x75)
value LANG_HEBREW (0x0d)
value LANG_HINDI (0x39)
value LANG_HUNGARIAN (0x0e)
value LANG_ICELANDIC (0x0f)
value LANG_IGBO (0x70)
value LANG_INDONESIAN (0x21)
value LANG_INUKTITUT (0x5d)
value LANG_INVARIANT (0x7f)
value LANG_IRISH (0x3c)
value LANG_ITALIAN (0x10)
value LANG_JAPANESE (0x11)
value LANG_KANNADA (0x4b)
value LANG_KASHMIRI (0x60)
value LANG_KAZAK (0x3f)
value LANG_KHMER (0x53)
value LANG_KICHE (0x86)
value LANG_KINYARWANDA (0x87)
value LANG_KONKANI (0x57)
value LANG_KOREAN (0x12)
value LANG_KYRGYZ (0x40)
value LANG_LAO (0x54)
value LANG_LATVIAN (0x26)
value LANG_LITHUANIAN (0x27)
value LANG_LOWER_SORBIAN (0x2e)
value LANG_LUXEMBOURGISH (0x6e)
value LANG_MACEDONIAN (0x2f)
value LANG_MALAY (0x3e)
value LANG_MALAYALAM (0x4c)
value LANG_MALTESE (0x3a)
value LANG_MANIPURI (0x58)
value LANG_MAORI (0x81)
value LANG_MAPUDUNGUN (0x7a)
value LANG_MARATHI (0x4e)
value LANG_MOHAWK (0x7c)
value LANG_MONGOLIAN (0x50)
value LANG_NEPALI (0x61)
value LANG_NEUTRAL (0x00)
value LANG_NORWEGIAN (0x14)
value LANG_OCCITAN (0x82)
value LANG_ODIA (0x48)
value LANG_ORIYA (0x48)
value LANG_PASHTO (0x63)
value LANG_PERSIAN (0x29)
value LANG_POLISH (0x15)
value LANG_PORTUGUESE (0x16)
value LANG_PULAR (0x67)
value LANG_PUNJABI (0x46)
value LANG_QUECHUA (0x6b)
value LANG_ROMANIAN (0x18)
value LANG_ROMANSH (0x17)
value LANG_RUSSIAN (0x19)
value LANG_SAKHA (0x85)
value LANG_SAMI (0x3b)
value LANG_SANSKRIT (0x4f)
value LANG_SCOTTISH_GAELIC (0x91)
value LANG_SERBIAN (0x1a)
value LANG_SERBIAN_NEUTRAL (0x7c1a)
value LANG_SINDHI (0x59)
value LANG_SINHALESE (0x5b)
value LANG_SLOVAK (0x1b)
value LANG_SLOVENIAN (0x24)
value LANG_SOTHO (0x6c)
value LANG_SPANISH (0x0a)
value LANG_SWAHILI (0x41)
value LANG_SWEDISH (0x1d)
value LANG_SYRIAC (0x5a)
value LANG_TAJIK (0x28)
value LANG_TAMAZIGHT (0x5f)
value LANG_TAMIL (0x49)
value LANG_TATAR (0x44)
value LANG_TELUGU (0x4a)
value LANG_THAI (0x1e)
value LANG_TIBETAN (0x51)
value LANG_TIGRIGNA (0x73)
value LANG_TIGRINYA (0x73)
value LANG_TSWANA (0x32)
value LANG_TURKISH (0x1f)
value LANG_TURKMEN (0x42)
value LANG_UIGHUR (0x80)
value LANG_UKRAINIAN (0x22)
value LANG_UPPER_SORBIAN (0x2e)
value LANG_URDU (0x20)
value LANG_UZBEK (0x43)
value LANG_VALENCIAN (0x03)
value LANG_VIETNAMESE (0x2a)
value LANG_WELSH (0x52)
value LANG_WOLOF (0x88)
value LANG_XHOSA (0x34)
value LANG_YAKUT (0x85)
value LANG_YI (0x78)
value LANG_YORUBA (0x6a)
value LANG_ZULU (0x35)
value LAYERED_PROTOCOL (0)
value LAYOUT_BITMAPORIENTATIONPRESERVED (0x00000008)
value LAYOUT_BTT (0x00000002)
value LAYOUT_ORIENTATIONMASK ((LAYOUT_RTL | LAYOUT_BTT | LAYOUT_VBH))
value LAYOUT_RTL (0x00000001)
value LAYOUT_VBH (0x00000004)
value LBN_DBLCLK (2)
value LBN_ERRSPACE ((-2))
value LBN_KILLFOCUS (5)
value LBN_SELCANCEL (3)
value LBN_SELCHANGE (1)
value LBN_SETFOCUS (4)
value LBSELCHSTRING (LBSELCHSTRINGA)
value LBS_COMBOBOX (0x8000L)
value LBS_DISABLENOSCROLL (0x1000L)
value LBS_EXTENDEDSEL (0x0800L)
value LBS_HASSTRINGS (0x0040L)
value LBS_MULTICOLUMN (0x0200L)
value LBS_MULTIPLESEL (0x0008L)
value LBS_NODATA (0x2000L)
value LBS_NOINTEGRALHEIGHT (0x0100L)
value LBS_NOREDRAW (0x0004L)
value LBS_NOSEL (0x4000L)
value LBS_NOTIFY (0x0001L)
value LBS_OWNERDRAWFIXED (0x0010L)
value LBS_OWNERDRAWVARIABLE (0x0020L)
value LBS_SORT (0x0002L)
value LBS_STANDARD ((LBS_NOTIFY | LBS_SORT | WS_VSCROLL | WS_BORDER))
value LBS_USETABSTOPS (0x0080L)
value LBS_WANTKEYBOARDINPUT (0x0400L)
value LB_ADDFILE (0x0196)
value LB_ADDSTRING (0x0180)
value LB_CTLCODE (0)
value LB_DELETESTRING (0x0182)
value LB_DIR (0x018D)
value LB_ERR ((-1))
value LB_ERRSPACE ((-2))
value LB_FINDSTRING (0x018F)
value LB_FINDSTRINGEXACT (0x01A2)
value LB_GETANCHORINDEX (0x019D)
value LB_GETCARETINDEX (0x019F)
value LB_GETCOUNT (0x018B)
value LB_GETCURSEL (0x0188)
value LB_GETHORIZONTALEXTENT (0x0193)
value LB_GETITEMDATA (0x0199)
value LB_GETITEMHEIGHT (0x01A1)
value LB_GETITEMRECT (0x0198)
value LB_GETLISTBOXINFO (0x01B2)
value LB_GETLOCALE (0x01A6)
value LB_GETSEL (0x0187)
value LB_GETSELCOUNT (0x0190)
value LB_GETSELITEMS (0x0191)
value LB_GETTEXT (0x0189)
value LB_GETTEXTLEN (0x018A)
value LB_GETTOPINDEX (0x018E)
value LB_INITSTORAGE (0x01A8)
value LB_INSERTSTRING (0x0181)
value LB_ITEMFROMPOINT (0x01A9)
value LB_MSGMAX (0x01B3)
value LB_OKAY (0)
value LB_RESETCONTENT (0x0184)
value LB_SELECTSTRING (0x018C)
value LB_SELITEMRANGE (0x019B)
value LB_SELITEMRANGEEX (0x0183)
value LB_SETANCHORINDEX (0x019C)
value LB_SETCARETINDEX (0x019E)
value LB_SETCOLUMNWIDTH (0x0195)
value LB_SETCOUNT (0x01A7)
value LB_SETCURSEL (0x0186)
value LB_SETHORIZONTALEXTENT (0x0194)
value LB_SETITEMDATA (0x019A)
value LB_SETITEMHEIGHT (0x01A0)
value LB_SETLOCALE (0x01A5)
value LB_SETSEL (0x0185)
value LB_SETTABSTOPS (0x0192)
value LB_SETTOPINDEX (0x0197)
value LCID_ALTERNATE_SORTS (0x00000004)
value LCID_INSTALLED (0x00000001)
value LCID_SUPPORTED (0x00000002)
value LCMAP_BYTEREV (0x00000800)
value LCMAP_FULLWIDTH (0x00800000)
value LCMAP_HALFWIDTH (0x00400000)
value LCMAP_HASH (0x00040000)
value LCMAP_HIRAGANA (0x00100000)
value LCMAP_KATAKANA (0x00200000)
value LCMAP_LINGUISTIC_CASING (0x01000000)
value LCMAP_LOWERCASE (0x00000100)
value LCMAP_SIMPLIFIED_CHINESE (0x02000000)
value LCMAP_SORTHANDLE (0x20000000)
value LCMAP_SORTKEY (0x00000400)
value LCMAP_TITLECASE (0x00000300)
value LCMAP_TRADITIONAL_CHINESE (0x04000000)
value LCMAP_UPPERCASE (0x00000200)
value LCS_CALIBRATED_RGB (0x00000000L)
value LCS_GM_ABS_COLORIMETRIC (0x00000008L)
value LCS_GM_BUSINESS (0x00000001L)
value LCS_GM_GRAPHICS (0x00000002L)
value LCS_GM_IMAGES (0x00000004L)
value LC_INTERIORS (128)
value LC_MARKER (4)
value LC_NONE (0)
value LC_POLYLINE (2)
value LC_POLYMARKER (8)
value LC_STYLED (32)
value LC_WIDE (16)
value LC_WIDESTYLED (64)
value LEFT_ALT_PRESSED (0x0002)
value LEFT_CTRL_PRESSED (0x0008)
value LF_FACESIZE (32)
value LF_FULLFACESIZE (64)
value LGRPID_ARABIC (0x000d)
value LGRPID_ARMENIAN (0x0011)
value LGRPID_BALTIC (0x0003)
value LGRPID_CENTRAL_EUROPE (0x0002)
value LGRPID_CYRILLIC (0x0005)
value LGRPID_GEORGIAN (0x0010)
value LGRPID_GREEK (0x0004)
value LGRPID_HEBREW (0x000c)
value LGRPID_INDIC (0x000f)
value LGRPID_INSTALLED (0x00000001)
value LGRPID_JAPANESE (0x0007)
value LGRPID_KOREAN (0x0008)
value LGRPID_SIMPLIFIED_CHINESE (0x000a)
value LGRPID_SUPPORTED (0x00000002)
value LGRPID_THAI (0x000b)
value LGRPID_TRADITIONAL_CHINESE (0x0009)
value LGRPID_TURKIC (0x0006)
value LGRPID_TURKISH (0x0006)
value LGRPID_VIETNAMESE (0x000e)
value LGRPID_WESTERN_EUROPE (0x0001)
value LHND ((LMEM_MOVEABLE | LMEM_ZEROINIT))
value LINECAPS (30)
value LINGUISTIC_IGNORECASE (0x00000010)
value LINGUISTIC_IGNOREDIACRITIC (0x00000020)
value LISTEN_OUTSTANDING (0x01)
value LITTLEENDIAN (0x0001)
value LLKHF_INJECTED (0x00000010)
value LLKHF_LOWER_IL_INJECTED (0x00000002)
value LLMHF_INJECTED (0x00000001)
value LLMHF_LOWER_IL_INJECTED (0x00000002)
value LMEM_DISCARDABLE (0x0F00)
value LMEM_DISCARDED (0x4000)
value LMEM_FIXED (0x0000)
value LMEM_INVALID_HANDLE (0x8000)
value LMEM_LOCKCOUNT (0x00FF)
value LMEM_MODIFY (0x0080)
value LMEM_MOVEABLE (0x0002)
value LMEM_NOCOMPACT (0x0010)
value LMEM_NODISCARD (0x0020)
value LMEM_VALID_FLAGS (0x0F72)
value LMEM_ZEROINIT (0x0040)
value LOAD_DLL_DEBUG_EVENT (6)
value LOAD_IGNORE_CODE_AUTHZ_LEVEL (0x00000010)
value LOAD_LIBRARY_AS_DATAFILE (0x00000002)
value LOAD_LIBRARY_AS_DATAFILE_EXCLUSIVE (0x00000040)
value LOAD_LIBRARY_AS_IMAGE_RESOURCE (0x00000020)
value LOAD_LIBRARY_OS_INTEGRITY_CONTINUITY (0x00008000)
value LOAD_LIBRARY_REQUIRE_SIGNED_TARGET (0x00000080)
value LOAD_LIBRARY_SAFE_CURRENT_DIRS (0x00002000)
value LOAD_LIBRARY_SEARCH_APPLICATION_DIR (0x00000200)
value LOAD_LIBRARY_SEARCH_DEFAULT_DIRS (0x00001000)
value LOAD_LIBRARY_SEARCH_DLL_LOAD_DIR (0x00000100)
value LOAD_LIBRARY_SEARCH_USER_DIRS (0x00000400)
value LOAD_WITH_ALTERED_SEARCH_PATH (0x00000008)
value LOCALE_ALL (0)
value LOCALE_ALLOW_NEUTRAL_NAMES (0x08000000)
value LOCALE_ALTERNATE_SORTS (0x00000004)
value LOCALE_ENUMPROC (LOCALE_ENUMPROCA)
value LOCALE_FONTSIGNATURE (0x00000058)
value LOCALE_ICALENDARTYPE (0x00001009)
value LOCALE_ICENTURY (0x00000024)
value LOCALE_ICONSTRUCTEDLOCALE (0x0000007d)
value LOCALE_ICOUNTRY (LOCALE_IDIALINGCODE)
value LOCALE_ICURRDIGITS (0x00000019)
value LOCALE_ICURRENCY (0x0000001B)
value LOCALE_IDATE (0x00000021)
value LOCALE_IDAYLZERO (0x00000026)
value LOCALE_IDEFAULTANSICODEPAGE (0x00001004)
value LOCALE_IDEFAULTCODEPAGE (0x0000000B)
value LOCALE_IDEFAULTCOUNTRY (0x0000000A)
value LOCALE_IDEFAULTEBCDICCODEPAGE (0x00001012)
value LOCALE_IDEFAULTLANGUAGE (0x00000009)
value LOCALE_IDEFAULTMACCODEPAGE (0x00001011)
value LOCALE_IDIALINGCODE (0x00000005)
value LOCALE_IDIGITS (0x00000011)
value LOCALE_IDIGITSUBSTITUTION (0x00001014)
value LOCALE_IFIRSTDAYOFWEEK (0x0000100C)
value LOCALE_IFIRSTWEEKOFYEAR (0x0000100D)
value LOCALE_IGEOID (0x0000005B)
value LOCALE_IINTLCURRDIGITS (0x0000001A)
value LOCALE_ILANGUAGE (0x00000001)
value LOCALE_ILDATE (0x00000022)
value LOCALE_ILZERO (0x00000012)
value LOCALE_IMEASURE (0x0000000D)
value LOCALE_IMONLZERO (0x00000027)
value LOCALE_INEGATIVEPERCENT (0x00000074)
value LOCALE_INEGCURR (0x0000001C)
value LOCALE_INEGNUMBER (0x00001010)
value LOCALE_INEGSEPBYSPACE (0x00000057)
value LOCALE_INEGSIGNPOSN (0x00000053)
value LOCALE_INEGSYMPRECEDES (0x00000056)
value LOCALE_INEUTRAL (0x00000071)
value LOCALE_IOPTIONALCALENDAR (0x0000100B)
value LOCALE_IPAPERSIZE (0x0000100A)
value LOCALE_IPOSITIVEPERCENT (0x00000075)
value LOCALE_IPOSSEPBYSPACE (0x00000055)
value LOCALE_IPOSSIGNPOSN (0x00000052)
value LOCALE_IPOSSYMPRECEDES (0x00000054)
value LOCALE_IREADINGLAYOUT (0x00000070)
value LOCALE_ITIME (0x00000023)
value LOCALE_ITIMEMARKPOSN (0x00001005)
value LOCALE_ITLZERO (0x00000025)
value LOCALE_NAME_MAX_LENGTH (85)
value LOCALE_NAME_USER_DEFAULT (NULL)
value LOCALE_NEUTRALDATA (0x00000010)
value LOCALE_NOUSEROVERRIDE (0x80000000)
value LOCALE_REPLACEMENT (0x00000008)
value LOCALE_RETURN_GENITIVE_NAMES (0x10000000)
value LOCALE_RETURN_NUMBER (0x20000000)
value LOCALE_SABBREVCTRYNAME (0x00000007)
value LOCALE_SABBREVLANGNAME (0x00000003)
value LOCALE_SAM (0x00000028)
value LOCALE_SCONSOLEFALLBACKNAME (0x0000006e)
value LOCALE_SCOUNTRY (LOCALE_SLOCALIZEDCOUNTRYNAME)
value LOCALE_SCURRENCY (0x00000014)
value LOCALE_SDATE (0x0000001D)
value LOCALE_SDECIMAL (0x0000000E)
value LOCALE_SDURATION (0x0000005d)
value LOCALE_SENGCOUNTRY (LOCALE_SENGLISHCOUNTRYNAME)
value LOCALE_SENGCURRNAME (0x00001007)
value LOCALE_SENGLANGUAGE (LOCALE_SENGLISHLANGUAGENAME)
value LOCALE_SENGLISHCOUNTRYNAME (0x00001002)
value LOCALE_SENGLISHDISPLAYNAME (0x00000072)
value LOCALE_SENGLISHLANGUAGENAME (0x00001001)
value LOCALE_SGROUPING (0x00000010)
value LOCALE_SINTLSYMBOL (0x00000015)
value LOCALE_SKEYBOARDSTOINSTALL (0x0000005e)
value LOCALE_SLANGDISPLAYNAME (LOCALE_SLOCALIZEDLANGUAGENAME)
value LOCALE_SLANGUAGE (LOCALE_SLOCALIZEDDISPLAYNAME)
value LOCALE_SLIST (0x0000000C)
value LOCALE_SLOCALIZEDCOUNTRYNAME (0x00000006)
value LOCALE_SLOCALIZEDDISPLAYNAME (0x00000002)
value LOCALE_SLOCALIZEDLANGUAGENAME (0x0000006f)
value LOCALE_SLONGDATE (0x00000020)
value LOCALE_SMONDECIMALSEP (0x00000016)
value LOCALE_SMONGROUPING (0x00000018)
value LOCALE_SMONTHDAY (0x00000078)
value LOCALE_SMONTHOUSANDSEP (0x00000017)
value LOCALE_SNAME (0x0000005c)
value LOCALE_SNAN (0x00000069)
value LOCALE_SNATIVECOUNTRYNAME (0x00000008)
value LOCALE_SNATIVECTRYNAME (LOCALE_SNATIVECOUNTRYNAME)
value LOCALE_SNATIVECURRNAME (0x00001008)
value LOCALE_SNATIVEDIGITS (0x00000013)
value LOCALE_SNATIVEDISPLAYNAME (0x00000073)
value LOCALE_SNATIVELANGNAME (LOCALE_SNATIVELANGUAGENAME)
value LOCALE_SNATIVELANGUAGENAME (0x00000004)
value LOCALE_SNEGATIVESIGN (0x00000051)
value LOCALE_SNEGINFINITY (0x0000006b)
value LOCALE_SOPENTYPELANGUAGETAG (0x0000007a)
value LOCALE_SPARENT (0x0000006d)
value LOCALE_SPECIFICDATA (0x00000020)
value LOCALE_SPERCENT (0x00000076)
value LOCALE_SPERMILLE (0x00000077)
value LOCALE_SPM (0x00000029)
value LOCALE_SPOSINFINITY (0x0000006a)
value LOCALE_SPOSITIVESIGN (0x00000050)
value LOCALE_SRELATIVELONGDATE (0x0000007c)
value LOCALE_SSCRIPTS (0x0000006c)
value LOCALE_SSHORTDATE (0x0000001F)
value LOCALE_SSHORTESTAM (0x0000007e)
value LOCALE_SSHORTESTPM (0x0000007f)
value LOCALE_SSHORTTIME (0x00000079)
value LOCALE_SSORTLOCALE (0x0000007b)
value LOCALE_SSORTNAME (0x00001013)
value LOCALE_STHOUSAND (0x0000000F)
value LOCALE_STIME (0x0000001E)
value LOCALE_STIMEFORMAT (0x00001003)
value LOCALE_SUPPLEMENTAL (0x00000002)
value LOCALE_SYEARMONTH (0x00001006)
value LOCALE_UNASSIGNED_LCID (LOCALE_CUSTOM_UNSPECIFIED)
value LOCALE_USE_CP_ACP (0x40000000)
value LOCALE_USE_NLS (0x10000000)
value LOCALE_WINDOWS (0x00000001)
value LOCKFILE_EXCLUSIVE_LOCK (0x00000002)
value LOCKFILE_FAIL_IMMEDIATELY (0x00000001)
value LOCK_ELEMENT (0)
value LOCK_UNLOCK_DOOR (0x02)
value LOCK_UNLOCK_IEPORT (0x01)
value LOCK_UNLOCK_KEYPAD (0x04)
value LOGON_NETCREDENTIALS_ONLY (0x00000002)
value LOGON_WITH_PROFILE (0x00000001)
value LOGON_ZERO_PASSWORD_BUFFER (0x80000000)
value LOGPIXELSX (88)
value LOGPIXELSY (90)
value LONG_MAX (2147483647)
value LONG_MIN ((-2147483647L - 1))
value LOOKUP_STREAM_FROM_CLUSTER_ENTRY_ATTRIBUTE_DATA (0x01000000)
value LOOKUP_STREAM_FROM_CLUSTER_ENTRY_ATTRIBUTE_INDEX (0x02000000)
value LOOKUP_STREAM_FROM_CLUSTER_ENTRY_ATTRIBUTE_MASK (0xff000000)
value LOOKUP_STREAM_FROM_CLUSTER_ENTRY_ATTRIBUTE_SYSTEM (0x03000000)
value LOOKUP_STREAM_FROM_CLUSTER_ENTRY_FLAG_DENY_DEFRAG_SET (0x00000002)
value LOOKUP_STREAM_FROM_CLUSTER_ENTRY_FLAG_FS_SYSTEM_FILE (0x00000004)
value LOOKUP_STREAM_FROM_CLUSTER_ENTRY_FLAG_PAGE_FILE (0x00000001)
value LOOKUP_STREAM_FROM_CLUSTER_ENTRY_FLAG_TXF_SYSTEM_FILE (0x00000008)
value LOW_SURROGATE_END (0xdfff)
value LOW_SURROGATE_START (0xdc00)
value LPCPROPSHEETHEADER (LPCPROPSHEETHEADERA)
value LPCPROPSHEETPAGE (LPCPROPSHEETPAGEA)
value LPCPROPSHEETPAGE_LATEST (LPCPROPSHEETPAGEA_LATEST)
value LPD_DOUBLEBUFFER (0x00000001)
value LPD_SHARE_ACCUM (0x00000100)
value LPD_SHARE_DEPTH (0x00000040)
value LPD_SHARE_STENCIL (0x00000080)
value LPD_STEREO (0x00000002)
value LPD_SUPPORT_GDI (0x00000010)
value LPD_SUPPORT_OPENGL (0x00000020)
value LPD_SWAP_COPY (0x00000400)
value LPD_SWAP_EXCHANGE (0x00000200)
value LPD_TRANSPARENT (0x00001000)
value LPD_TYPE_COLORINDEX (1)
value LPD_TYPE_RGBA (0)
value LPFNPSPCALLBACK (LPFNPSPCALLBACKA)
value LPOCNCONNPROC (LPOCNCONNPROCA)
value LPOINET (LPIINTERNET)
value LPOINETBINDINFO (LPIINTERNETBINDINFO)
value LPOINETPRIORITY (LPIINTERNETPRIORITY)
value LPOINETPROTOCOL (LPIINTERNETPROTOCOL)
value LPOINETPROTOCOLEX (LPIINTERNETPROTOCOLEX)
value LPOINETPROTOCOLINFO (LPIINTERNETPROTOCOLINFO)
value LPOINETPROTOCOLROOT (LPIINTERNETPROTOCOLROOT)
value LPOINETPROTOCOLSINK (LPIINTERNETPROTOCOLSINK)
value LPOINETPROTOCOLSINKSTACKABLE (LPIINTERNETPROTOCOLSINKSTACKABLE)
value LPOINETSESSION (LPIINTERNETSESSION)
value LPOINETTHREADSWITCH (LPIINTERNETTHREADSWITCH)
value LPOPENCARDNAMEA_EX (LPOPENCARDNAME_EXA)
value LPOPENCARDNAMEW_EX (LPOPENCARDNAME_EXW)
value LPOPENCARDNAME_A (LPOPENCARDNAMEA)
value LPOPENCARDNAME_W (LPOPENCARDNAMEW)
value LPPROPSHEETHEADER (LPPROPSHEETHEADERA)
value LPPROPSHEETPAGE (LPPROPSHEETPAGEA)
value LPPROPSHEETPAGE_LATEST (LPPROPSHEETPAGEA_LATEST)
value LPSCARD_READERSTATE_A (LPSCARD_READERSTATEA)
value LPSCARD_READERSTATE_W (LPSCARD_READERSTATEW)
value LPSERVICE_MAIN_FUNCTION (LPSERVICE_MAIN_FUNCTIONA)
value LPTR ((LMEM_FIXED | LMEM_ZEROINIT))
value LPWSAEVENT (LPHANDLE)
value LR_COLOR (0x00000002)
value LR_COPYDELETEORG (0x00000008)
value LR_COPYFROMRESOURCE (0x00004000)
value LR_COPYRETURNORG (0x00000004)
value LR_CREATEDIBSECTION (0x00002000)
value LR_DEFAULTCOLOR (0x00000000)
value LR_DEFAULTSIZE (0x00000040)
value LR_LOADFROMFILE (0x00000010)
value LR_LOADTRANSPARENT (0x00000020)
value LR_MONOCHROME (0x00000001)
value LR_SHARED (0x00008000)
value LR_VGACOLOR (0x00000080)
value LSFW_LOCK (1)
value LSFW_UNLOCK (2)
value LTGRAY_BRUSH (1)
value LTP_PC_SMT (0x1)
value LUA_TOKEN (0x4)
value LUP_ADDRCONFIG (0x00100000)
value LUP_API_ANSI (0x01000000)
value LUP_CONTAINERS (0x00000002)
value LUP_DEEP (0x00000001)
value LUP_DISABLE_IDN_ENCODING (0x00800000)
value LUP_DNS_ONLY (0x00020000)
value LUP_DUAL_ADDR (0x00200000)
value LUP_EXCLUSIVE_CUSTOM_SERVERS (0x08000000)
value LUP_EXTENDED_QUERYSET (0x02000000)
value LUP_FILESERVER (0x00400000)
value LUP_FLUSHCACHE (0x00001000)
value LUP_FLUSHPREVIOUS (0x00002000)
value LUP_FORCE_CLEAR_TEXT (0x40000000)
value LUP_NEAREST (0x00000008)
value LUP_NOCONTAINERS (0x00000004)
value LUP_NON_AUTHORITATIVE (0x00004000)
value LUP_REQUIRE_SECURE (0x10000000)
value LUP_RESOLUTION_HANDLE (0x80000000)
value LUP_RES_SERVICE (0x00008000)
value LUP_RETURN_ADDR (0x00000100)
value LUP_RETURN_ALIASES (0x00000400)
value LUP_RETURN_ALL (0x00000FF0)
value LUP_RETURN_BLOB (0x00000200)
value LUP_RETURN_COMMENT (0x00000080)
value LUP_RETURN_NAME (0x00000010)
value LUP_RETURN_PREFERRED_NAMES (0x00010000)
value LUP_RETURN_QUERY_STRING (0x00000800)
value LUP_RETURN_RESPONSE_FLAGS (0x00040000)
value LUP_RETURN_TTL (0x20000000)
value LUP_RETURN_TYPE (0x00000020)
value LUP_RETURN_VERSION (0x00000040)
value LUP_SECURE (0x00008000)
value LUP_SECURE_WITH_FALLBACK (0x04000000)
value LWA_ALPHA (0x00000002)
value LWA_COLORKEY (0x00000001)
value LZERROR_BADINHANDLE ((-1))
value LZERROR_BADOUTHANDLE ((-2))
value LZERROR_BADVALUE ((-7))
value LZERROR_GLOBALLOC ((-5))
value LZERROR_GLOBLOCK ((-6))
value LZERROR_READ ((-3))
value LZERROR_UNKNOWNALG ((-8))
value LZERROR_WRITE ((-4))
value MAC_CHARSET (77)
value MAILSLOT_NO_MESSAGE (((DWORD)-1))
value MAILSLOT_WAIT_FOREVER (((DWORD)-1))
value MAKEINTRESOURCE (MAKEINTRESOURCEA)
value MAPVK_VK_TO_CHAR ((2))
value MAPVK_VK_TO_VSC ((0))
value MAPVK_VK_TO_VSC_EX ((4))
value MAPVK_VSC_TO_VK ((1))
value MAPVK_VSC_TO_VK_EX ((3))
value MAP_COMPOSITE (0x00000040)
value MAP_EXPAND_LIGATURES (0x00002000)
value MAP_FOLDCZONE (0x00000010)
value MAP_FOLDDIGITS (0x00000080)
value MAP_PRECOMPOSED (0x00000020)
value MARKPARITY (3)
value MARK_HANDLE_CLOUD_SYNC ((0x00000800))
value MARK_HANDLE_DISABLE_FILE_METADATA_OPTIMIZATION ((0x00001000))
value MARK_HANDLE_ENABLE_CPU_CACHE ((0x10000000))
value MARK_HANDLE_ENABLE_USN_SOURCE_ON_PAGING_IO ((0x00002000))
value MARK_HANDLE_FILTER_METADATA ((0x00000200))
value MARK_HANDLE_NOT_READ_COPY ((0x00000100))
value MARK_HANDLE_NOT_REALTIME ((0x00000040))
value MARK_HANDLE_NOT_TXF_SYSTEM_LOG ((0x00000008))
value MARK_HANDLE_PROTECT_CLUSTERS ((0x00000001))
value MARK_HANDLE_READ_COPY ((0x00000080))
value MARK_HANDLE_REALTIME ((0x00000020))
value MARK_HANDLE_RETURN_PURGE_FAILURE ((0x00000400))
value MARK_HANDLE_SKIP_COHERENCY_SYNC_DISALLOW_WRITES ((0x00004000))
value MARK_HANDLE_SUPPRESS_VOLUME_OPEN_FLUSH ((0x00008000))
value MARK_HANDLE_TXF_SYSTEM_LOG ((0x00000004))
value MARSHALINTERFACE_MIN (500)
value MARSHAL_E_FIRST (0x80040120L)
value MARSHAL_E_LAST (0x8004012FL)
value MARSHAL_S_FIRST (0x00040120L)
value MARSHAL_S_LAST (0x0004012FL)
value MAXBYTE (0xff)
value MAXCHAR (0x7f)
value MAXDWORD (0xffffffff)
value MAXERRORLENGTH (256)
value MAXGETHOSTSTRUCT (1024)
value MAXIMUM_ALLOWED ((0x02000000L))
value MAXIMUM_ATTR_STRING_LENGTH (32)
value MAXIMUM_ENCRYPTION_VALUE (0x00000004)
value MAXIMUM_PROCESSORS (MAXIMUM_PROC_PER_GROUP)
value MAXIMUM_PROC_PER_GROUP (64)
value MAXIMUM_RESERVED_MANIFEST_RESOURCE_ID (MAKEINTRESOURCE(16 ))
value MAXIMUM_SMARTCARD_READERS (10)
value MAXIMUM_SUSPEND_COUNT (MAXCHAR)
value MAXIMUM_WAIT_OBJECTS (64)
value MAXIMUM_XSTATE_FEATURES ((64))
value MAXINTATOM (0xC000)
value MAXLOGICALLOGNAMESIZE (256)
value MAXLONG (0x7fffffff)
value MAXPNAMELEN (32)
value MAXPROPPAGES (100)
value MAXSHORT (0x7fff)
value MAXSTRETCHBLTMODE (4)
value MAXUIDLEN (64)
value MAXWORD (0xffff)
value MAX_ACL_REVISION (ACL_REVISION4)
value MAX_COMPUTERNAME_LENGTH (15)
value MAX_DEFAULTCHAR (2)
value MAX_FORM_KEYWORD_LENGTH (63+1)
value MAX_FW_BUCKET_ID_LENGTH (132)
value MAX_HW_COUNTERS (16)
value MAX_INTERFACE_CODES (8)
value MAX_JOYSTICKOEMVXDNAME (260)
value MAX_LANA (254)
value MAX_LEADBYTES (12)
value MAX_LOGICALDPIOVERRIDE (2)
value MAX_MONITORS (4)
value MAX_NUM_REASONS (256)
value MAX_PATH (260)
value MAX_PERF_OBJECTS_IN_QUERY_FUNCTION ((64L))
value MAX_PRIORITY (99)
value MAX_PROFILE_LEN (80)
value MAX_PROTOCOL_CHAIN (7)
value MAX_REASON_BUGID_LEN (32)
value MAX_REASON_COMMENT_LEN (512)
value MAX_REASON_DESC_LEN (256)
value MAX_REASON_NAME_LEN (64)
value MAX_RESOURCEMANAGER_DESCRIPTION_LENGTH (64)
value MAX_SID_SIZE (256)
value MAX_SIZE_SECURITY_ID (512)
value MAX_STR_BLOCKREASON (256)
value MAX_TOUCH_COUNT (256)
value MAX_TOUCH_PREDICTION_FILTER_TAPS (3)
value MAX_TRANSACTION_DESCRIPTION_LENGTH (64)
value MAX_UCSCHAR ((0x0010FFFF))
value MAX_VOLUME_ID_SIZE (36)
value MAX_VOLUME_TEMPLATE_SIZE (40)
value MA_ACTIVATE (1)
value MA_ACTIVATEANDEAT (2)
value MA_NOACTIVATE (3)
value MA_NOACTIVATEANDEAT (4)
value MB_ABORTRETRYIGNORE (0x00000002L)
value MB_APPLMODAL (0x00000000L)
value MB_CANCELTRYCONTINUE (0x00000006L)
value MB_COMPOSITE (0x00000002)
value MB_DEFAULT_DESKTOP_ONLY (0x00020000L)
value MB_DEFMASK (0x00000F00L)
value MB_ERR_INVALID_CHARS (0x00000008)
value MB_HELP (0x00004000L)
value MB_ICONASTERISK (0x00000040L)
value MB_ICONERROR (MB_ICONHAND)
value MB_ICONEXCLAMATION (0x00000030L)
value MB_ICONHAND (0x00000010L)
value MB_ICONINFORMATION (MB_ICONASTERISK)
value MB_ICONMASK (0x000000F0L)
value MB_ICONQUESTION (0x00000020L)
value MB_ICONSTOP (MB_ICONHAND)
value MB_ICONWARNING (MB_ICONEXCLAMATION)
value MB_LEN_MAX (5)
value MB_MISCMASK (0x0000C000L)
value MB_MODEMASK (0x00003000L)
value MB_NOFOCUS (0x00008000L)
value MB_OK (0x00000000L)
value MB_OKCANCEL (0x00000001L)
value MB_PRECOMPOSED (0x00000001)
value MB_RETRYCANCEL (0x00000005L)
value MB_RIGHT (0x00080000L)
value MB_RTLREADING (0x00100000L)
value MB_SERVICE_NOTIFICATION (0x00200000L)
value MB_SETFOREGROUND (0x00010000L)
value MB_SYSTEMMODAL (0x00001000L)
value MB_TASKMODAL (0x00002000L)
value MB_TOPMOST (0x00040000L)
value MB_TYPEMASK (0x0000000FL)
value MB_USEGLYPHCHARS (0x00000004)
value MB_USERICON (0x00000080L)
value MB_YESNO (0x00000004L)
value MB_YESNOCANCEL (0x00000003L)
value MCIERR_BAD_CONSTANT ((MCIERR_BASE + 34))
value MCIERR_BAD_INTEGER ((MCIERR_BASE + 14))
value MCIERR_BAD_TIME_FORMAT ((MCIERR_BASE + 37))
value MCIERR_BASE (256)
value MCIERR_CANNOT_LOAD_DRIVER ((MCIERR_BASE + 10))
value MCIERR_CANNOT_USE_ALL ((MCIERR_BASE + 23))
value MCIERR_CREATEWINDOW ((MCIERR_BASE + 91))
value MCIERR_CUSTOM_DRIVER_BASE ((MCIERR_BASE + 256))
value MCIERR_DEVICE_LENGTH ((MCIERR_BASE + 54))
value MCIERR_DEVICE_LOCKED ((MCIERR_BASE + 32))
value MCIERR_DEVICE_NOT_INSTALLED ((MCIERR_BASE + 50))
value MCIERR_DEVICE_NOT_READY ((MCIERR_BASE + 20))
value MCIERR_DEVICE_OPEN ((MCIERR_BASE + 9))
value MCIERR_DEVICE_ORD_LENGTH ((MCIERR_BASE + 55))
value MCIERR_DEVICE_TYPE_REQUIRED ((MCIERR_BASE + 31))
value MCIERR_DRIVER ((MCIERR_BASE + 22))
value MCIERR_DRIVER_INTERNAL ((MCIERR_BASE + 16))
value MCIERR_DUPLICATE_ALIAS ((MCIERR_BASE + 33))
value MCIERR_DUPLICATE_FLAGS ((MCIERR_BASE + 39))
value MCIERR_EXTENSION_NOT_FOUND ((MCIERR_BASE + 25))
value MCIERR_EXTRA_CHARACTERS ((MCIERR_BASE + 49))
value MCIERR_FILENAME_REQUIRED ((MCIERR_BASE + 48))
value MCIERR_FILE_NOT_FOUND ((MCIERR_BASE + 19))
value MCIERR_FILE_NOT_SAVED ((MCIERR_BASE + 30))
value MCIERR_FILE_READ ((MCIERR_BASE + 92))
value MCIERR_FILE_WRITE ((MCIERR_BASE + 93))
value MCIERR_FLAGS_NOT_COMPATIBLE ((MCIERR_BASE + 28))
value MCIERR_GET_CD ((MCIERR_BASE + 51))
value MCIERR_HARDWARE ((MCIERR_BASE + 6))
value MCIERR_ILLEGAL_FOR_AUTO_OPEN ((MCIERR_BASE + 47))
value MCIERR_INTERNAL ((MCIERR_BASE + 21))
value MCIERR_INVALID_DEVICE_ID ((MCIERR_BASE + 1))
value MCIERR_INVALID_DEVICE_NAME ((MCIERR_BASE + 7))
value MCIERR_INVALID_FILE ((MCIERR_BASE + 40))
value MCIERR_MISSING_COMMAND_STRING ((MCIERR_BASE + 11))
value MCIERR_MISSING_DEVICE_NAME ((MCIERR_BASE + 36))
value MCIERR_MISSING_PARAMETER ((MCIERR_BASE + 17))
value MCIERR_MISSING_STRING_ARGUMENT ((MCIERR_BASE + 13))
value MCIERR_MULTIPLE ((MCIERR_BASE + 24))
value MCIERR_MUST_USE_SHAREABLE ((MCIERR_BASE + 35))
value MCIERR_NEW_REQUIRES_ALIAS ((MCIERR_BASE + 43))
value MCIERR_NONAPPLICABLE_FUNCTION ((MCIERR_BASE + 46))
value MCIERR_NOTIFY_ON_AUTO_OPEN ((MCIERR_BASE + 44))
value MCIERR_NO_CLOSING_QUOTE ((MCIERR_BASE + 38))
value MCIERR_NO_ELEMENT_ALLOWED ((MCIERR_BASE + 45))
value MCIERR_NO_IDENTITY ((MCIERR_BASE + 94))
value MCIERR_NO_INTEGER ((MCIERR_BASE + 56))
value MCIERR_NO_WINDOW ((MCIERR_BASE + 90))
value MCIERR_NULL_PARAMETER_BLOCK ((MCIERR_BASE + 41))
value MCIERR_OUTOFRANGE ((MCIERR_BASE + 26))
value MCIERR_OUT_OF_MEMORY ((MCIERR_BASE + 8))
value MCIERR_PARAM_OVERFLOW ((MCIERR_BASE + 12))
value MCIERR_PARSER_INTERNAL ((MCIERR_BASE + 15))
value MCIERR_SEQ_DIV_INCOMPATIBLE ((MCIERR_BASE + 80))
value MCIERR_SEQ_NOMIDIPRESENT ((MCIERR_BASE + 87))
value MCIERR_SEQ_PORTUNSPECIFIED ((MCIERR_BASE + 86))
value MCIERR_SEQ_PORT_INUSE ((MCIERR_BASE + 81))
value MCIERR_SEQ_PORT_MAPNODEVICE ((MCIERR_BASE + 83))
value MCIERR_SEQ_PORT_MISCERROR ((MCIERR_BASE + 84))
value MCIERR_SEQ_PORT_NONEXISTENT ((MCIERR_BASE + 82))
value MCIERR_SEQ_TIMER ((MCIERR_BASE + 85))
value MCIERR_SET_CD ((MCIERR_BASE + 52))
value MCIERR_SET_DRIVE ((MCIERR_BASE + 53))
value MCIERR_UNNAMED_RESOURCE ((MCIERR_BASE + 42))
value MCIERR_UNRECOGNIZED_COMMAND ((MCIERR_BASE + 5))
value MCIERR_UNRECOGNIZED_KEYWORD ((MCIERR_BASE + 3))
value MCIERR_UNSUPPORTED_FUNCTION ((MCIERR_BASE + 18))
value MCIERR_WAVE_INPUTSINUSE ((MCIERR_BASE + 66))
value MCIERR_WAVE_INPUTSUNSUITABLE ((MCIERR_BASE + 72))
value MCIERR_WAVE_INPUTUNSPECIFIED ((MCIERR_BASE + 69))
value MCIERR_WAVE_OUTPUTSINUSE ((MCIERR_BASE + 64))
value MCIERR_WAVE_OUTPUTSUNSUITABLE ((MCIERR_BASE + 70))
value MCIERR_WAVE_OUTPUTUNSPECIFIED ((MCIERR_BASE + 68))
value MCIERR_WAVE_SETINPUTINUSE ((MCIERR_BASE + 67))
value MCIERR_WAVE_SETINPUTUNSUITABLE ((MCIERR_BASE + 73))
value MCIERR_WAVE_SETOUTPUTINUSE ((MCIERR_BASE + 65))
value MCIERR_WAVE_SETOUTPUTUNSUITABLE ((MCIERR_BASE + 71))
value MCI_ALL_DEVICE_ID (((MCIDEVICEID)-1))
value MCI_ANIM_GETDEVCAPS_CAN_REVERSE (0x00004001L)
value MCI_ANIM_GETDEVCAPS_CAN_STRETCH (0x00004007L)
value MCI_ANIM_GETDEVCAPS_FAST_RATE (0x00004002L)
value MCI_ANIM_GETDEVCAPS_MAX_WINDOWS (0x00004008L)
value MCI_ANIM_GETDEVCAPS_NORMAL_RATE (0x00004004L)
value MCI_ANIM_GETDEVCAPS_PALETTES (0x00004006L)
value MCI_ANIM_GETDEVCAPS_SLOW_RATE (0x00004003L)
value MCI_ANIM_INFO_TEXT (0x00010000L)
value MCI_ANIM_OPEN_NOSTATIC (0x00040000L)
value MCI_ANIM_OPEN_PARENT (0x00020000L)
value MCI_ANIM_OPEN_WS (0x00010000L)
value MCI_ANIM_PLAY_FAST (0x00040000L)
value MCI_ANIM_PLAY_REVERSE (0x00020000L)
value MCI_ANIM_PLAY_SCAN (0x00100000L)
value MCI_ANIM_PLAY_SLOW (0x00080000L)
value MCI_ANIM_PLAY_SPEED (0x00010000L)
value MCI_ANIM_PUT_DESTINATION (0x00040000L)
value MCI_ANIM_PUT_SOURCE (0x00020000L)
value MCI_ANIM_REALIZE_BKGD (0x00020000L)
value MCI_ANIM_REALIZE_NORM (0x00010000L)
value MCI_ANIM_RECT (0x00010000L)
value MCI_ANIM_STATUS_FORWARD (0x00004002L)
value MCI_ANIM_STATUS_HPAL (0x00004004L)
value MCI_ANIM_STATUS_HWND (0x00004003L)
value MCI_ANIM_STATUS_SPEED (0x00004001L)
value MCI_ANIM_STATUS_STRETCH (0x00004005L)
value MCI_ANIM_STEP_FRAMES (0x00020000L)
value MCI_ANIM_STEP_REVERSE (0x00010000L)
value MCI_ANIM_UPDATE_HDC (0x00020000L)
value MCI_ANIM_WHERE_DESTINATION (0x00040000L)
value MCI_ANIM_WHERE_SOURCE (0x00020000L)
value MCI_ANIM_WINDOW_DEFAULT (0x00000000L)
value MCI_ANIM_WINDOW_DISABLE_STRETCH (0x00200000L)
value MCI_ANIM_WINDOW_ENABLE_STRETCH (0x00100000L)
value MCI_ANIM_WINDOW_HWND (0x00010000L)
value MCI_ANIM_WINDOW_STATE (0x00040000L)
value MCI_ANIM_WINDOW_TEXT (0x00080000L)
value MCI_BREAK (0x0811)
value MCI_BREAK_HWND (0x00000200L)
value MCI_BREAK_KEY (0x00000100L)
value MCI_BREAK_OFF (0x00000400L)
value MCI_CDA_STATUS_TYPE_TRACK (0x00004001L)
value MCI_CDA_TRACK_AUDIO ((MCI_CD_OFFSET + 0))
value MCI_CDA_TRACK_OTHER ((MCI_CD_OFFSET + 1))
value MCI_CD_OFFSET (1088)
value MCI_CLOSE (0x0804)
value MCI_COPY (0x0852)
value MCI_CUE (0x0830)
value MCI_CUT (0x0851)
value MCI_DELETE (0x0856)
value MCI_DEVTYPE_ANIMATION (519)
value MCI_DEVTYPE_CD_AUDIO (516)
value MCI_DEVTYPE_DAT (517)
value MCI_DEVTYPE_DIGITAL_VIDEO (520)
value MCI_DEVTYPE_FIRST (MCI_DEVTYPE_VCR)
value MCI_DEVTYPE_FIRST_USER (0x1000)
value MCI_DEVTYPE_LAST (MCI_DEVTYPE_SEQUENCER)
value MCI_DEVTYPE_OTHER (521)
value MCI_DEVTYPE_OVERLAY (515)
value MCI_DEVTYPE_SCANNER (518)
value MCI_DEVTYPE_SEQUENCER (523)
value MCI_DEVTYPE_VCR (513)
value MCI_DEVTYPE_VIDEODISC (514)
value MCI_DEVTYPE_WAVEFORM_AUDIO (522)
value MCI_ESCAPE (0x0805)
value MCI_FIRST (DRV_MCI_FIRST)
value MCI_FORMAT_BYTES (8)
value MCI_FORMAT_FRAMES (3)
value MCI_FORMAT_HMS (1)
value MCI_FORMAT_MILLISECONDS (0)
value MCI_FORMAT_MSF (2)
value MCI_FORMAT_SAMPLES (9)
value MCI_FORMAT_TMSF (10)
value MCI_FREEZE (0x0844)
value MCI_FROM (0x00000004L)
value MCI_GETDEVCAPS (0x080B)
value MCI_GETDEVCAPS_CAN_EJECT (0x00000007L)
value MCI_GETDEVCAPS_CAN_PLAY (0x00000008L)
value MCI_GETDEVCAPS_CAN_RECORD (0x00000001L)
value MCI_GETDEVCAPS_CAN_SAVE (0x00000009L)
value MCI_GETDEVCAPS_COMPOUND_DEVICE (0x00000006L)
value MCI_GETDEVCAPS_DEVICE_TYPE (0x00000004L)
value MCI_GETDEVCAPS_HAS_AUDIO (0x00000002L)
value MCI_GETDEVCAPS_HAS_VIDEO (0x00000003L)
value MCI_GETDEVCAPS_ITEM (0x00000100L)
value MCI_GETDEVCAPS_USES_FILES (0x00000005L)
value MCI_INFO (0x080A)
value MCI_INFO_COPYRIGHT (0x00002000L)
value MCI_INFO_FILE (0x00000200L)
value MCI_INFO_MEDIA_IDENTITY (0x00000800L)
value MCI_INFO_MEDIA_UPC (0x00000400L)
value MCI_INFO_NAME (0x00001000L)
value MCI_INFO_PRODUCT (0x00000100L)
value MCI_LAST (0x0FFF)
value MCI_LOAD (0x0850)
value MCI_LOAD_FILE (0x00000100L)
value MCI_MODE_NOT_READY ((MCI_STRING_OFFSET + 12))
value MCI_MODE_OPEN ((MCI_STRING_OFFSET + 18))
value MCI_MODE_PAUSE ((MCI_STRING_OFFSET + 17))
value MCI_MODE_PLAY ((MCI_STRING_OFFSET + 14))
value MCI_MODE_RECORD ((MCI_STRING_OFFSET + 15))
value MCI_MODE_SEEK ((MCI_STRING_OFFSET + 16))
value MCI_MODE_STOP ((MCI_STRING_OFFSET + 13))
value MCI_NOTIFY (0x00000001L)
value MCI_NOTIFY_ABORTED (0x0004)
value MCI_NOTIFY_FAILURE (0x0008)
value MCI_NOTIFY_SUCCESSFUL (0x0001)
value MCI_NOTIFY_SUPERSEDED (0x0002)
value MCI_OPEN (0x0803)
value MCI_OPEN_ALIAS (0x00000400L)
value MCI_OPEN_ELEMENT (0x00000200L)
value MCI_OPEN_ELEMENT_ID (0x00000800L)
value MCI_OPEN_SHAREABLE (0x00000100L)
value MCI_OPEN_TYPE (0x00002000L)
value MCI_OPEN_TYPE_ID (0x00001000L)
value MCI_OVLY_GETDEVCAPS_CAN_FREEZE (0x00004002L)
value MCI_OVLY_GETDEVCAPS_CAN_STRETCH (0x00004001L)
value MCI_OVLY_GETDEVCAPS_MAX_WINDOWS (0x00004003L)
value MCI_OVLY_INFO_TEXT (0x00010000L)
value MCI_OVLY_OPEN_PARENT (0x00020000L)
value MCI_OVLY_OPEN_WS (0x00010000L)
value MCI_OVLY_PUT_DESTINATION (0x00040000L)
value MCI_OVLY_PUT_FRAME (0x00080000L)
value MCI_OVLY_PUT_SOURCE (0x00020000L)
value MCI_OVLY_PUT_VIDEO (0x00100000L)
value MCI_OVLY_RECT (0x00010000L)
value MCI_OVLY_STATUS_HWND (0x00004001L)
value MCI_OVLY_STATUS_STRETCH (0x00004002L)
value MCI_OVLY_WHERE_DESTINATION (0x00040000L)
value MCI_OVLY_WHERE_FRAME (0x00080000L)
value MCI_OVLY_WHERE_SOURCE (0x00020000L)
value MCI_OVLY_WHERE_VIDEO (0x00100000L)
value MCI_OVLY_WINDOW_DEFAULT (0x00000000L)
value MCI_OVLY_WINDOW_DISABLE_STRETCH (0x00200000L)
value MCI_OVLY_WINDOW_ENABLE_STRETCH (0x00100000L)
value MCI_OVLY_WINDOW_HWND (0x00010000L)
value MCI_OVLY_WINDOW_STATE (0x00040000L)
value MCI_OVLY_WINDOW_TEXT (0x00080000L)
value MCI_PASTE (0x0853)
value MCI_PAUSE (0x0809)
value MCI_PLAY (0x0806)
value MCI_PUT (0x0842)
value MCI_REALIZE (0x0840)
value MCI_RECORD (0x080F)
value MCI_RECORD_INSERT (0x00000100L)
value MCI_RECORD_OVERWRITE (0x00000200L)
value MCI_RESUME (0x0855)
value MCI_SAVE (0x0813)
value MCI_SAVE_FILE (0x00000100L)
value MCI_SEEK (0x0807)
value MCI_SEEK_TO_END (0x00000200L)
value MCI_SEEK_TO_START (0x00000100L)
value MCI_SEQ_DIV_PPQN ((0 + MCI_SEQ_OFFSET))
value MCI_SEQ_FILE (0x4002)
value MCI_SEQ_FORMAT_SONGPTR (0x4001)
value MCI_SEQ_MAPPER (65535)
value MCI_SEQ_MIDI (0x4003)
value MCI_SEQ_NONE (65533)
value MCI_SEQ_OFFSET (1216)
value MCI_SEQ_SET_MASTER (0x00080000L)
value MCI_SEQ_SET_OFFSET (0x01000000L)
value MCI_SEQ_SET_PORT (0x00020000L)
value MCI_SEQ_SET_SLAVE (0x00040000L)
value MCI_SEQ_SET_TEMPO (0x00010000L)
value MCI_SEQ_SMPTE (0x4004)
value MCI_SEQ_STATUS_COPYRIGHT (0x0000400CL)
value MCI_SEQ_STATUS_DIVTYPE (0x0000400AL)
value MCI_SEQ_STATUS_MASTER (0x00004008L)
value MCI_SEQ_STATUS_NAME (0x0000400BL)
value MCI_SEQ_STATUS_OFFSET (0x00004009L)
value MCI_SEQ_STATUS_PORT (0x00004003L)
value MCI_SEQ_STATUS_SLAVE (0x00004007L)
value MCI_SEQ_STATUS_TEMPO (0x00004002L)
value MCI_SET (0x080D)
value MCI_SET_AUDIO (0x00000800L)
value MCI_SET_AUDIO_ALL (0x00000000L)
value MCI_SET_AUDIO_LEFT (0x00000001L)
value MCI_SET_AUDIO_RIGHT (0x00000002L)
value MCI_SET_DOOR_CLOSED (0x00000200L)
value MCI_SET_DOOR_OPEN (0x00000100L)
value MCI_SET_OFF (0x00004000L)
value MCI_SET_ON (0x00002000L)
value MCI_SET_TIME_FORMAT (0x00000400L)
value MCI_SET_VIDEO (0x00001000L)
value MCI_SPIN (0x080C)
value MCI_STATUS (0x0814)
value MCI_STATUS_CURRENT_TRACK (0x00000008L)
value MCI_STATUS_ITEM (0x00000100L)
value MCI_STATUS_LENGTH (0x00000001L)
value MCI_STATUS_MEDIA_PRESENT (0x00000005L)
value MCI_STATUS_MODE (0x00000004L)
value MCI_STATUS_NUMBER_OF_TRACKS (0x00000003L)
value MCI_STATUS_POSITION (0x00000002L)
value MCI_STATUS_READY (0x00000007L)
value MCI_STATUS_START (0x00000200L)
value MCI_STATUS_TIME_FORMAT (0x00000006L)
value MCI_STEP (0x080E)
value MCI_STOP (0x0808)
value MCI_STRING_OFFSET (512)
value MCI_SYSINFO (0x0810)
value MCI_SYSINFO_INSTALLNAME (0x00000800L)
value MCI_SYSINFO_NAME (0x00000400L)
value MCI_SYSINFO_OPEN (0x00000200L)
value MCI_SYSINFO_QUANTITY (0x00000100L)
value MCI_TO (0x00000008L)
value MCI_TRACK (0x00000010L)
value MCI_UNFREEZE (0x0845)
value MCI_UPDATE (0x0854)
value MCI_USER_MESSAGES ((DRV_MCI_FIRST + 0x400))
value MCI_VD_ESCAPE_STRING (0x00000100L)
value MCI_VD_FORMAT_TRACK (0x4001)
value MCI_VD_GETDEVCAPS_CAN_REVERSE (0x00004002L)
value MCI_VD_GETDEVCAPS_CAV (0x00020000L)
value MCI_VD_GETDEVCAPS_CLV (0x00010000L)
value MCI_VD_GETDEVCAPS_FAST_RATE (0x00004003L)
value MCI_VD_GETDEVCAPS_NORMAL_RATE (0x00004005L)
value MCI_VD_GETDEVCAPS_SLOW_RATE (0x00004004L)
value MCI_VD_MEDIA_CAV ((MCI_VD_OFFSET + 3))
value MCI_VD_MEDIA_CLV ((MCI_VD_OFFSET + 2))
value MCI_VD_MEDIA_OTHER ((MCI_VD_OFFSET + 4))
value MCI_VD_MODE_PARK ((MCI_VD_OFFSET + 1))
value MCI_VD_OFFSET (1024)
value MCI_VD_PLAY_FAST (0x00020000L)
value MCI_VD_PLAY_REVERSE (0x00010000L)
value MCI_VD_PLAY_SCAN (0x00080000L)
value MCI_VD_PLAY_SLOW (0x00100000L)
value MCI_VD_PLAY_SPEED (0x00040000L)
value MCI_VD_SEEK_REVERSE (0x00010000L)
value MCI_VD_SPIN_DOWN (0x00020000L)
value MCI_VD_SPIN_UP (0x00010000L)
value MCI_VD_STATUS_DISC_SIZE (0x00004006L)
value MCI_VD_STATUS_FORWARD (0x00004003L)
value MCI_VD_STATUS_MEDIA_TYPE (0x00004004L)
value MCI_VD_STATUS_SIDE (0x00004005L)
value MCI_VD_STATUS_SPEED (0x00004002L)
value MCI_VD_STEP_FRAMES (0x00010000L)
value MCI_VD_STEP_REVERSE (0x00020000L)
value MCI_WAIT (0x00000002L)
value MCI_WAVE_GETDEVCAPS_INPUTS (0x00004001L)
value MCI_WAVE_GETDEVCAPS_OUTPUTS (0x00004002L)
value MCI_WAVE_INPUT (0x00400000L)
value MCI_WAVE_MAPPER ((MCI_WAVE_OFFSET + 1))
value MCI_WAVE_OFFSET (1152)
value MCI_WAVE_OPEN_BUFFER (0x00010000L)
value MCI_WAVE_OUTPUT (0x00800000L)
value MCI_WAVE_PCM ((MCI_WAVE_OFFSET + 0))
value MCI_WAVE_SET_ANYINPUT (0x04000000L)
value MCI_WAVE_SET_ANYOUTPUT (0x08000000L)
value MCI_WAVE_SET_AVGBYTESPERSEC (0x00080000L)
value MCI_WAVE_SET_BITSPERSAMPLE (0x00200000L)
value MCI_WAVE_SET_BLOCKALIGN (0x00100000L)
value MCI_WAVE_SET_CHANNELS (0x00020000L)
value MCI_WAVE_SET_FORMATTAG (0x00010000L)
value MCI_WAVE_SET_SAMPLESPERSEC (0x00040000L)
value MCI_WAVE_STATUS_AVGBYTESPERSEC (0x00004004L)
value MCI_WAVE_STATUS_BITSPERSAMPLE (0x00004006L)
value MCI_WAVE_STATUS_BLOCKALIGN (0x00004005L)
value MCI_WAVE_STATUS_CHANNELS (0x00004002L)
value MCI_WAVE_STATUS_FORMATTAG (0x00004001L)
value MCI_WAVE_STATUS_LEVEL (0x00004007L)
value MCI_WAVE_STATUS_SAMPLESPERSEC (0x00004003L)
value MCI_WHERE (0x0843)
value MCI_WINDOW (0x0841)
value MDIS_ALLCHILDSTYLES (0x0001)
value MDITILE_HORIZONTAL (0x0001)
value MDITILE_SKIPDISABLED (0x0002)
value MDITILE_VERTICAL (0x0000)
value MDITILE_ZORDER (0x0004)
value MDMSPKRFLAG_CALLSETUP (0x00000008)
value MDMSPKRFLAG_DIAL (0x00000002)
value MDMSPKRFLAG_OFF (0x00000001)
value MDMSPKRFLAG_ON (0x00000004)
value MDMSPKR_CALLSETUP (0x00000003)
value MDMSPKR_DIAL (0x00000001)
value MDMSPKR_OFF (0x00000000)
value MDMSPKR_ON (0x00000002)
value MDMVOLFLAG_HIGH (0x00000004)
value MDMVOLFLAG_LOW (0x00000001)
value MDMVOLFLAG_MEDIUM (0x00000002)
value MDMVOL_HIGH (0x00000002)
value MDMVOL_LOW (0x00000000)
value MDMVOL_MEDIUM (0x00000001)
value MDM_ANALOG_RLP_OFF (0x1)
value MDM_ANALOG_RLP_ON (0x0)
value MDM_AUTO_ML_DEFAULT (0x0)
value MDM_AUTO_ML_NONE (0x1)
value MDM_AUTO_SPEED_DEFAULT (0x0)
value MDM_BEARERMODE_ANALOG (0x0)
value MDM_BEARERMODE_GSM (0x2)
value MDM_BEARERMODE_ISDN (0x1)
value MDM_BLIND_DIAL (0x00000200)
value MDM_CCITT_OVERRIDE (0x00000040)
value MDM_CELLULAR (0x00000008)
value MDM_COMPRESSION (0x00000001)
value MDM_DIAGNOSTICS (0x00000800)
value MDM_ERROR_CONTROL (0x00000002)
value MDM_FLOWCONTROL_HARD (0x00000010)
value MDM_FLOWCONTROL_SOFT (0x00000020)
value MDM_FORCED_EC (0x00000004)
value MDM_HDLCPPP_AUTH_CHAP (0x3)
value MDM_HDLCPPP_AUTH_DEFAULT (0x0)
value MDM_HDLCPPP_AUTH_MSCHAP (0x4)
value MDM_HDLCPPP_AUTH_NONE (0x1)
value MDM_HDLCPPP_AUTH_PAP (0x2)
value MDM_HDLCPPP_ML_DEFAULT (0x0)
value MDM_HDLCPPP_ML_NONE (0x1)
value MDM_HDLCPPP_SPEED_DEFAULT (0x0)
value MDM_MASK_AUTO_SPEED (0x7)
value MDM_MASK_BEARERMODE (0x0000f000)
value MDM_MASK_EXTENDEDINFO ((MDM_MASK_BEARERMODE|MDM_MASK_PROTOCOLINFO))
value MDM_MASK_HDLCPPP_SPEED (0x7)
value MDM_MASK_PROTOCOLDATA (0x0ff00000)
value MDM_MASK_PROTOCOLID (0x000f0000)
value MDM_MASK_PROTOCOLINFO ((MDM_MASK_PROTOCOLID|MDM_MASK_PROTOCOLDATA))
value MDM_PIAFS_INCOMING (0)
value MDM_PIAFS_OUTGOING (1)
value MDM_PROTOCOLID_ANALOG (0x7)
value MDM_PROTOCOLID_AUTO (0x6)
value MDM_PROTOCOLID_DEFAULT (0x0)
value MDM_PROTOCOLID_GPRS (0x8)
value MDM_PROTOCOLID_HDLCPPP (0x1)
value MDM_PROTOCOLID_PIAFS (0x9)
value MDM_SHIFT_AUTO_ML (0x6)
value MDM_SHIFT_AUTO_SPEED (0x0)
value MDM_SHIFT_BEARERMODE (12)
value MDM_SHIFT_EXTENDEDINFO (MDM_SHIFT_BEARERMODE)
value MDM_SHIFT_HDLCPPP_AUTH (0x3)
value MDM_SHIFT_HDLCPPP_ML (0x6)
value MDM_SHIFT_HDLCPPP_SPEED (0x0)
value MDM_SHIFT_PROTOCOLDATA (20)
value MDM_SHIFT_PROTOCOLID (16)
value MDM_SHIFT_PROTOCOLINFO (MDM_SHIFT_PROTOCOLID)
value MDM_SPEED_ADJUST (0x00000080)
value MDM_TONE_DIAL (0x00000100)
value MEDIA_CURRENTLY_MOUNTED (0x80000000)
value MEDIA_ERASEABLE (0x00000001)
value MEDIA_READ_ONLY (0x00000004)
value MEDIA_READ_WRITE (0x00000008)
value MEDIA_WRITE_ONCE (0x00000002)
value MEDIA_WRITE_PROTECTED (0x00000100)
value MEHC_PATROL_SCRUBBER_PRESENT (0x1)
value MEMBERID_NIL (DISPID_UNKNOWN)
value MEMORY_ALLOCATION_ALIGNMENT (16)
value MEMORY_CURRENT_PARTITION_HANDLE (((HANDLE) (LONG_PTR) -1))
value MEMORY_EXISTING_VAD_PARTITION_HANDLE (((HANDLE) (LONG_PTR) -3))
value MEMORY_PARTITION_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | SYNCHRONIZE | MEMORY_PARTITION_QUERY_ACCESS | MEMORY_PARTITION_MODIFY_ACCESS))
value MEMORY_PARTITION_MODIFY_ACCESS (0x0002)
value MEMORY_PARTITION_QUERY_ACCESS (0x0001)
value MEMORY_PRIORITY_BELOW_NORMAL (4)
value MEMORY_PRIORITY_LOW (2)
value MEMORY_PRIORITY_LOWEST (0)
value MEMORY_PRIORITY_MEDIUM (3)
value MEMORY_PRIORITY_NORMAL (5)
value MEMORY_PRIORITY_VERY_LOW (1)
value MEMORY_SYSTEM_PARTITION_HANDLE (((HANDLE) (LONG_PTR) -2))
value MEM_COALESCE_PLACEHOLDERS (0x00000001)
value MEM_COMMIT (0x00001000)
value MEM_DECOMMIT (0x00004000)
value MEM_DEDICATED_ATTRIBUTE_NOT_SPECIFIED (((DWORD64) -1))
value MEM_DIFFERENT_IMAGE_BASE_OK (0x00800000)
value MEM_EXTENDED_PARAMETER_EC_CODE (0x00000040)
value MEM_EXTENDED_PARAMETER_GRAPHICS (0x00000001)
value MEM_EXTENDED_PARAMETER_IMAGE_NO_HPAT (0x00000080)
value MEM_EXTENDED_PARAMETER_NONPAGED (0x00000002)
value MEM_EXTENDED_PARAMETER_NONPAGED_HUGE (0x00000010)
value MEM_EXTENDED_PARAMETER_NONPAGED_LARGE (0x00000008)
value MEM_EXTENDED_PARAMETER_NUMA_NODE_MANDATORY (MINLONG64)
value MEM_EXTENDED_PARAMETER_SOFT_FAULT_PAGES (0x00000020)
value MEM_EXTENDED_PARAMETER_TYPE_BITS (8)
value MEM_EXTENDED_PARAMETER_ZERO_PAGES_OPTIONAL (0x00000004)
value MEM_E_INVALID_LINK (_HRESULT_TYPEDEF_(0x80080010L))
value MEM_E_INVALID_ROOT (_HRESULT_TYPEDEF_(0x80080009L))
value MEM_E_INVALID_SIZE (_HRESULT_TYPEDEF_(0x80080011L))
value MEM_FREE (0x00010000)
value MEM_IMAGE (0x01000000)
value MEM_LARGE_PAGES (0x20000000)
value MEM_MAPPED (0x00040000)
value MEM_PHYSICAL (0x00400000)
value MEM_PRESERVE_PLACEHOLDER (0x00000002)
value MEM_PRIVATE (0x00020000)
value MEM_RELEASE (0x00008000)
value MEM_REPLACE_PLACEHOLDER (0x00004000)
value MEM_RESERVE (0x00002000)
value MEM_RESERVE_PLACEHOLDER (0x00040000)
value MEM_RESET (0x00080000)
value MEM_RESET_UNDO (0x01000000)
value MEM_ROTATE (0x00800000)
value MEM_TOP_DOWN (0x00100000)
value MEM_UNMAP_WITH_TRANSIENT_BOOST (0x00000001)
value MEM_WRITE_WATCH (0x00200000)
value MENROLL_E_CERTAUTH_FAILED_TO_FIND_CERT (_HRESULT_TYPEDEF_(0x80180028L))
value MENROLL_E_CERTPOLICY_PRIVATEKEYCREATION_FAILED (_HRESULT_TYPEDEF_(0x80180027L))
value MENROLL_E_CONNECTIVITY (_HRESULT_TYPEDEF_(0x80180010L))
value MENROLL_E_DEVICECAPREACHED (_HRESULT_TYPEDEF_(0x80180013L))
value MENROLL_E_DEVICENOTSUPPORTED (_HRESULT_TYPEDEF_(0x80180014L))
value MENROLL_E_DEVICE_ALREADY_ENROLLED (_HRESULT_TYPEDEF_(0x8018000AL))
value MENROLL_E_DEVICE_AUTHENTICATION_ERROR (_HRESULT_TYPEDEF_(0x80180002L))
value MENROLL_E_DEVICE_AUTHORIZATION_ERROR (_HRESULT_TYPEDEF_(0x80180003L))
value MENROLL_E_DEVICE_CERTIFICATEREQUEST_ERROR (_HRESULT_TYPEDEF_(0x80180004L))
value MENROLL_E_DEVICE_CONFIGMGRSERVER_ERROR (_HRESULT_TYPEDEF_(0x80180005L))
value MENROLL_E_DEVICE_INTERNALSERVICE_ERROR (_HRESULT_TYPEDEF_(0x80180006L))
value MENROLL_E_DEVICE_INVALIDSECURITY_ERROR (_HRESULT_TYPEDEF_(0x80180007L))
value MENROLL_E_DEVICE_MANAGEMENT_BLOCKED (_HRESULT_TYPEDEF_(0x80180026L))
value MENROLL_E_DEVICE_MESSAGE_FORMAT_ERROR (_HRESULT_TYPEDEF_(0x80180001L))
value MENROLL_E_DEVICE_UNKNOWN_ERROR (_HRESULT_TYPEDEF_(0x80180008L))
value MENROLL_E_DISCOVERY_SEC_CERT_DATE_INVALID (_HRESULT_TYPEDEF_(0x8018000DL))
value MENROLL_E_EMPTY_MESSAGE (_HRESULT_TYPEDEF_(0x80180029L))
value MENROLL_E_ENROLLMENTDATAINVALID (_HRESULT_TYPEDEF_(0x80180019L))
value MENROLL_E_ENROLLMENT_IN_PROGRESS (_HRESULT_TYPEDEF_(0x80180009L))
value MENROLL_E_INMAINTENANCE (_HRESULT_TYPEDEF_(0x80180017L))
value MENROLL_E_INSECUREREDIRECT (_HRESULT_TYPEDEF_(0x8018001AL))
value MENROLL_E_INVALIDSSLCERT (_HRESULT_TYPEDEF_(0x80180012L))
value MENROLL_E_MDM_NOT_CONFIGURED (_HRESULT_TYPEDEF_(0x80180031L))
value MENROLL_E_NOTELIGIBLETORENEW (_HRESULT_TYPEDEF_(0x80180016L))
value MENROLL_E_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80180015L))
value MENROLL_E_PASSWORD_NEEDED (_HRESULT_TYPEDEF_(0x8018000EL))
value MENROLL_E_PLATFORM_LICENSE_ERROR (_HRESULT_TYPEDEF_(0x8018001CL))
value MENROLL_E_PLATFORM_UNKNOWN_ERROR (_HRESULT_TYPEDEF_(0x8018001DL))
value MENROLL_E_PLATFORM_WRONG_STATE (_HRESULT_TYPEDEF_(0x8018001BL))
value MENROLL_E_PROV_CSP_APPMGMT (_HRESULT_TYPEDEF_(0x80180025L))
value MENROLL_E_PROV_CSP_CERTSTORE (_HRESULT_TYPEDEF_(0x8018001EL))
value MENROLL_E_PROV_CSP_DMCLIENT (_HRESULT_TYPEDEF_(0x80180020L))
value MENROLL_E_PROV_CSP_MISC (_HRESULT_TYPEDEF_(0x80180022L))
value MENROLL_E_PROV_CSP_PFW (_HRESULT_TYPEDEF_(0x80180021L))
value MENROLL_E_PROV_SSLCERTNOTFOUND (_HRESULT_TYPEDEF_(0x80180024L))
value MENROLL_E_PROV_UNKNOWN (_HRESULT_TYPEDEF_(0x80180023L))
value MENROLL_E_USER_CANCELLED (_HRESULT_TYPEDEF_(0x80180030L))
value MENROLL_E_USER_LICENSE (_HRESULT_TYPEDEF_(0x80180018L))
value MENROLL_E_WAB_ERROR (_HRESULT_TYPEDEF_(0x8018000FL))
value MENROLL_S_ENROLLMENT_SUSPENDED (_HRESULT_TYPEDEF_(0x00180011L))
value MENU_EVENT (0x0008)
value MERGECOPY ((DWORD)0x00C000CA)
value MERGEPAINT ((DWORD)0x00BB0226)
value MESSAGE_RESOURCE_UNICODE (0x0001)
value METAFILE_DRIVER (2049)
value META_ANIMATEPALETTE (0x0436)
value META_ARC (0x0817)
value META_BITBLT (0x0922)
value META_CHORD (0x0830)
value META_CREATEBRUSHINDIRECT (0x02FC)
value META_CREATEFONTINDIRECT (0x02FB)
value META_CREATEPALETTE (0x00f7)
value META_CREATEPATTERNBRUSH (0x01F9)
value META_CREATEPENINDIRECT (0x02FA)
value META_CREATEREGION (0x06FF)
value META_DELETEOBJECT (0x01f0)
value META_DIBBITBLT (0x0940)
value META_DIBCREATEPATTERNBRUSH (0x0142)
value META_DIBSTRETCHBLT (0x0b41)
value META_ELLIPSE (0x0418)
value META_ESCAPE (0x0626)
value META_EXCLUDECLIPRECT (0x0415)
value META_EXTFLOODFILL (0x0548)
value META_EXTTEXTOUT (0x0a32)
value META_FILLREGION (0x0228)
value META_FLOODFILL (0x0419)
value META_FRAMEREGION (0x0429)
value META_INTERSECTCLIPRECT (0x0416)
value META_INVERTREGION (0x012A)
value META_LINETO (0x0213)
value META_MOVETO (0x0214)
value META_OFFSETCLIPRGN (0x0220)
value META_OFFSETVIEWPORTORG (0x0211)
value META_OFFSETWINDOWORG (0x020F)
value META_PAINTREGION (0x012B)
value META_PATBLT (0x061D)
value META_PIE (0x081A)
value META_POLYGON (0x0324)
value META_POLYLINE (0x0325)
value META_POLYPOLYGON (0x0538)
value META_REALIZEPALETTE (0x0035)
value META_RECTANGLE (0x041B)
value META_RESIZEPALETTE (0x0139)
value META_RESTOREDC (0x0127)
value META_ROUNDRECT (0x061C)
value META_SAVEDC (0x001E)
value META_SCALEVIEWPORTEXT (0x0412)
value META_SCALEWINDOWEXT (0x0410)
value META_SELECTCLIPREGION (0x012C)
value META_SELECTOBJECT (0x012D)
value META_SELECTPALETTE (0x0234)
value META_SETBKCOLOR (0x0201)
value META_SETBKMODE (0x0102)
value META_SETDIBTODEV (0x0d33)
value META_SETLAYOUT (0x0149)
value META_SETMAPMODE (0x0103)
value META_SETMAPPERFLAGS (0x0231)
value META_SETPALENTRIES (0x0037)
value META_SETPIXEL (0x041F)
value META_SETPOLYFILLMODE (0x0106)
value META_SETRELABS (0x0105)
value META_SETSTRETCHBLTMODE (0x0107)
value META_SETTEXTALIGN (0x012E)
value META_SETTEXTCHAREXTRA (0x0108)
value META_SETTEXTCOLOR (0x0209)
value META_SETTEXTJUSTIFICATION (0x020A)
value META_SETVIEWPORTEXT (0x020E)
value META_SETVIEWPORTORG (0x020D)
value META_SETWINDOWEXT (0x020C)
value META_SETWINDOWORG (0x020B)
value META_STRETCHBLT (0x0B23)
value META_STRETCHDIB (0x0f43)
value META_TEXTOUT (0x0521)
value METHOD_BUFFERED (0)
value METHOD_DIRECT_FROM_HARDWARE (METHOD_OUT_DIRECT)
value METHOD_DIRECT_TO_HARDWARE (METHOD_IN_DIRECT)
value METHOD_IN_DIRECT (1)
value METHOD_NEITHER (3)
value METHOD_OUT_DIRECT (2)
value METRICS_USEDEFAULT (-1)
value MEVT_COMMENT (((BYTE)0x82))
value MEVT_F_CALLBACK (0x40000000L)
value MEVT_F_LONG (0x80000000L)
value MEVT_F_SHORT (0x00000000L)
value MEVT_LONGMSG (((BYTE)0x80))
value MEVT_NOP (((BYTE)0x02))
value MEVT_SHORTMSG (((BYTE)0x00))
value MEVT_TEMPO (((BYTE)0x01))
value MEVT_VERSION (((BYTE)0x84))
value MFCOMMENT (15)
value MFS_CHECKED (MF_CHECKED)
value MFS_DEFAULT (MF_DEFAULT)
value MFS_DISABLED (MFS_GRAYED)
value MFS_ENABLED (MF_ENABLED)
value MFS_GRAYED (0x00000003L)
value MFS_HILITE (MF_HILITE)
value MFS_UNCHECKED (MF_UNCHECKED)
value MFS_UNHILITE (MF_UNHILITE)
value MFT_BITMAP (MF_BITMAP)
value MFT_MENUBARBREAK (MF_MENUBARBREAK)
value MFT_MENUBREAK (MF_MENUBREAK)
value MFT_OWNERDRAW (MF_OWNERDRAW)
value MFT_RADIOCHECK (0x00000200L)
value MFT_RIGHTJUSTIFY (MF_RIGHTJUSTIFY)
value MFT_RIGHTORDER (0x00002000L)
value MFT_SEPARATOR (MF_SEPARATOR)
value MFT_STRING (MF_STRING)
value MF_APPEND (0x00000100L)
value MF_BITMAP (0x00000004L)
value MF_BYCOMMAND (0x00000000L)
value MF_BYPOSITION (0x00000400L)
value MF_CALLBACKS (0x08000000)
value MF_CHANGE (0x00000080L)
value MF_CHECKED (0x00000008L)
value MF_CONV (0x40000000)
value MF_DEFAULT (0x00001000L)
value MF_DELETE (0x00000200L)
value MF_DISABLED (0x00000002L)
value MF_ENABLED (0x00000000L)
value MF_END (0x00000080L)
value MF_ERRORS (0x10000000)
value MF_GRAYED (0x00000001L)
value MF_HELP (0x00004000L)
value MF_HILITE (0x00000080L)
value MF_HSZ_INFO (0x01000000)
value MF_INSERT (0x00000000L)
value MF_LINKS (0x20000000)
value MF_MASK (0xFF000000)
value MF_MENUBARBREAK (0x00000020L)
value MF_MENUBREAK (0x00000040L)
value MF_MOUSESELECT (0x00008000L)
value MF_OWNERDRAW (0x00000100L)
value MF_POPUP (0x00000010L)
value MF_POSTMSGS (0x04000000)
value MF_REMOVE (0x00001000L)
value MF_RIGHTJUSTIFY (0x00004000L)
value MF_SENDMSGS (0x02000000)
value MF_SEPARATOR (0x00000800L)
value MF_STRING (0x00000000L)
value MF_SYSMENU (0x00002000L)
value MF_UNCHECKED (0x00000000L)
value MF_UNHILITE (0x00000000L)
value MF_USECHECKBITMAPS (0x00000200L)
value MHDR_DONE (0x00000001)
value MHDR_INQUEUE (0x00000004)
value MHDR_ISSTRM (0x00000008)
value MHDR_PREPARED (0x00000002)
value MH_CLEANUP (4)
value MH_CREATE (1)
value MH_DELETE (3)
value MH_KEEP (2)
value MICROSOFT_ROOT_CERT_CHAIN_POLICY_CHECK_APPLICATION_ROOT_FLAG (0x00020000)
value MICROSOFT_ROOT_CERT_CHAIN_POLICY_DISABLE_FLIGHT_ROOT_FLAG (0x00040000)
value MICROSOFT_ROOT_CERT_CHAIN_POLICY_ENABLE_TEST_ROOT_FLAG (0x00010000)
value MICROSOFT_WINBASE_H_DEFINE_INTERLOCKED_CPLUSPLUS_OVERLOADS (0)
value MICROSOFT_WINDOWS_WINBASE_H_DEFINE_INTERLOCKED_CPLUSPLUS_OVERLOADS (1)
value MIDICAPS_CACHE (0x0004)
value MIDICAPS_LRVOLUME (0x0002)
value MIDICAPS_STREAM (0x0008)
value MIDICAPS_VOLUME (0x0001)
value MIDIERR_BADOPENMODE ((MIDIERR_BASE + 6))
value MIDIERR_BASE (64)
value MIDIERR_DONT_CONTINUE ((MIDIERR_BASE + 7))
value MIDIERR_INVALIDSETUP ((MIDIERR_BASE + 5))
value MIDIERR_LASTERROR ((MIDIERR_BASE + 7))
value MIDIERR_NODEVICE ((MIDIERR_BASE + 4))
value MIDIERR_NOMAP ((MIDIERR_BASE + 2))
value MIDIERR_NOTREADY ((MIDIERR_BASE + 3))
value MIDIERR_STILLPLAYING ((MIDIERR_BASE + 1))
value MIDIERR_UNPREPARED ((MIDIERR_BASE + 0))
value MIDIMAPPER (((UINT)-1))
value MIDIPATCHSIZE (128)
value MIDIPROP_GET (0x40000000L)
value MIDIPROP_SET (0x80000000L)
value MIDIPROP_TEMPO (0x00000002L)
value MIDIPROP_TIMEDIV (0x00000001L)
value MIDISTRM_ERROR ((-2))
value MIDI_CACHE_ALL (1)
value MIDI_CACHE_BESTFIT (2)
value MIDI_CACHE_QUERY (3)
value MIDI_IO_STATUS (0x00000020L)
value MIDI_MAPPER (((UINT)-1))
value MIDI_UNCACHE (4)
value MIIM_BITMAP (0x00000080)
value MIIM_CHECKMARKS (0x00000008)
value MIIM_DATA (0x00000020)
value MIIM_FTYPE (0x00000100)
value MIIM_ID (0x00000002)
value MIIM_STATE (0x00000001)
value MIIM_STRING (0x00000040)
value MIIM_SUBMENU (0x00000004)
value MIIM_TYPE (0x00000010)
value MILAVERR_INSUFFICIENTVIDEORESOURCES (_HRESULT_TYPEDEF_(0x88980508L))
value MILAVERR_INVALIDWMPVERSION (_HRESULT_TYPEDEF_(0x88980507L))
value MILAVERR_MEDIAPLAYERCLOSED (_HRESULT_TYPEDEF_(0x8898050DL))
value MILAVERR_MODULENOTLOADED (_HRESULT_TYPEDEF_(0x88980505L))
value MILAVERR_NOCLOCK (_HRESULT_TYPEDEF_(0x88980500L))
value MILAVERR_NOMEDIATYPE (_HRESULT_TYPEDEF_(0x88980501L))
value MILAVERR_NOREADYFRAMES (_HRESULT_TYPEDEF_(0x88980504L))
value MILAVERR_NOVIDEOMIXER (_HRESULT_TYPEDEF_(0x88980502L))
value MILAVERR_NOVIDEOPRESENTER (_HRESULT_TYPEDEF_(0x88980503L))
value MILAVERR_REQUESTEDTEXTURETOOBIG (_HRESULT_TYPEDEF_(0x8898050AL))
value MILAVERR_SEEKFAILED (_HRESULT_TYPEDEF_(0x8898050BL))
value MILAVERR_UNEXPECTEDWMPFAILURE (_HRESULT_TYPEDEF_(0x8898050CL))
value MILAVERR_UNKNOWNHARDWAREERROR (_HRESULT_TYPEDEF_(0x8898050EL))
value MILAVERR_VIDEOACCELERATIONNOTAVAILABLE (_HRESULT_TYPEDEF_(0x88980509L))
value MILAVERR_WMPFACTORYNOTREGISTERED (_HRESULT_TYPEDEF_(0x88980506L))
value MILCORE_TS_QUERYVER_RESULT_FALSE (0x0)
value MILCORE_TS_QUERYVER_RESULT_TRUE (0x7FFFFFFF)
value MILEFFECTSERR_ALREADYATTACHEDTOLISTENER (_HRESULT_TYPEDEF_(0x88980618L))
value MILEFFECTSERR_CONNECTORNOTASSOCIATEDWITHEFFECT (_HRESULT_TYPEDEF_(0x88980612L))
value MILEFFECTSERR_CONNECTORNOTCONNECTED (_HRESULT_TYPEDEF_(0x88980611L))
value MILEFFECTSERR_CYCLEDETECTED (_HRESULT_TYPEDEF_(0x88980614L))
value MILEFFECTSERR_EFFECTALREADYINAGRAPH (_HRESULT_TYPEDEF_(0x88980616L))
value MILEFFECTSERR_EFFECTHASNOCHILDREN (_HRESULT_TYPEDEF_(0x88980617L))
value MILEFFECTSERR_EFFECTINMORETHANONEGRAPH (_HRESULT_TYPEDEF_(0x88980615L))
value MILEFFECTSERR_EFFECTNOTPARTOFGROUP (_HRESULT_TYPEDEF_(0x8898060FL))
value MILEFFECTSERR_EMPTYBOUNDS (_HRESULT_TYPEDEF_(0x8898061AL))
value MILEFFECTSERR_NOINPUTSOURCEATTACHED (_HRESULT_TYPEDEF_(0x88980610L))
value MILEFFECTSERR_NOTAFFINETRANSFORM (_HRESULT_TYPEDEF_(0x88980619L))
value MILEFFECTSERR_OUTPUTSIZETOOLARGE (_HRESULT_TYPEDEF_(0x8898061BL))
value MILEFFECTSERR_RESERVED (_HRESULT_TYPEDEF_(0x88980613L))
value MILEFFECTSERR_UNKNOWNPROPERTY (_HRESULT_TYPEDEF_(0x8898060EL))
value MILERR_ADAPTER_NOT_FOUND (_HRESULT_TYPEDEF_(0x8898009EL))
value MILERR_ALREADYLOCKED (_HRESULT_TYPEDEF_(0x88980086L))
value MILERR_ALREADY_INITIALIZED (_HRESULT_TYPEDEF_(0x8898008FL))
value MILERR_BADNUMBER (_HRESULT_TYPEDEF_(0x8898000AL))
value MILERR_COLORSPACE_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8898009FL))
value MILERR_DEVICECANNOTRENDERTEXT (_HRESULT_TYPEDEF_(0x88980088L))
value MILERR_DISPLAYFORMATNOTSUPPORTED (_HRESULT_TYPEDEF_(0x88980084L))
value MILERR_DISPLAYID_ACCESS_DENIED (_HRESULT_TYPEDEF_(0x889800A1L))
value MILERR_DISPLAYSTATEINVALID (_HRESULT_TYPEDEF_(0x88980006L))
value MILERR_DXGI_ENUMERATION_OUT_OF_SYNC (_HRESULT_TYPEDEF_(0x8898009DL))
value MILERR_GENERIC_IGNORE (_HRESULT_TYPEDEF_(0x8898008BL))
value MILERR_GLYPHBITMAPMISSED (_HRESULT_TYPEDEF_(0x88980089L))
value MILERR_INSUFFICIENTBUFFER (_HRESULT_TYPEDEF_(0x88980002L))
value MILERR_INTERNALERROR (_HRESULT_TYPEDEF_(0x88980080L))
value MILERR_INVALIDCALL (_HRESULT_TYPEDEF_(0x88980085L))
value MILERR_MALFORMEDGLYPHCACHE (_HRESULT_TYPEDEF_(0x8898008AL))
value MILERR_MALFORMED_GUIDELINE_DATA (_HRESULT_TYPEDEF_(0x8898008CL))
value MILERR_MAX_TEXTURE_SIZE_EXCEEDED (_HRESULT_TYPEDEF_(0x8898009AL))
value MILERR_MISMATCHED_SIZE (_HRESULT_TYPEDEF_(0x88980090L))
value MILERR_MROW_READLOCK_FAILED (_HRESULT_TYPEDEF_(0x88980097L))
value MILERR_MROW_UPDATE_FAILED (_HRESULT_TYPEDEF_(0x88980098L))
value MILERR_NEED_RECREATE_AND_PRESENT (_HRESULT_TYPEDEF_(0x8898008EL))
value MILERR_NONINVERTIBLEMATRIX (_HRESULT_TYPEDEF_(0x88980007L))
value MILERR_NOTLOCKED (_HRESULT_TYPEDEF_(0x88980087L))
value MILERR_NOT_QUEUING_PRESENTS (_HRESULT_TYPEDEF_(0x88980094L))
value MILERR_NO_HARDWARE_DEVICE (_HRESULT_TYPEDEF_(0x8898008DL))
value MILERR_NO_REDIRECTION_SURFACE_AVAILABLE (_HRESULT_TYPEDEF_(0x88980091L))
value MILERR_NO_REDIRECTION_SURFACE_RETRY_LATER (_HRESULT_TYPEDEF_(0x88980095L))
value MILERR_OBJECTBUSY (_HRESULT_TYPEDEF_(0x88980001L))
value MILERR_PREFILTER_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x889800A0L))
value MILERR_QPC_TIME_WENT_BACKWARD (_HRESULT_TYPEDEF_(0x8898009BL))
value MILERR_QUEUED_PRESENT_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x88980093L))
value MILERR_REMOTING_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x88980092L))
value MILERR_SCANNER_FAILED (_HRESULT_TYPEDEF_(0x88980004L))
value MILERR_SCREENACCESSDENIED (_HRESULT_TYPEDEF_(0x88980005L))
value MILERR_SHADER_COMPILE_FAILED (_HRESULT_TYPEDEF_(0x88980099L))
value MILERR_TERMINATED (_HRESULT_TYPEDEF_(0x88980009L))
value MILERR_TOOMANYSHADERELEMNTS (_HRESULT_TYPEDEF_(0x88980096L))
value MILERR_ZEROVECTOR (_HRESULT_TYPEDEF_(0x88980008L))
value MIM_APPLYTOSUBMENUS (0x80000000)
value MIM_BACKGROUND (0x00000002)
value MIM_CLOSE (MM_MIM_CLOSE)
value MIM_DATA (MM_MIM_DATA)
value MIM_ERROR (MM_MIM_ERROR)
value MIM_HELPID (0x00000004)
value MIM_LONGDATA (MM_MIM_LONGDATA)
value MIM_LONGERROR (MM_MIM_LONGERROR)
value MIM_MAXHEIGHT (0x00000001)
value MIM_MENUDATA (0x00000008)
value MIM_MOREDATA (MM_MIM_MOREDATA)
value MIM_OPEN (MM_MIM_OPEN)
value MIM_STYLE (0x00000010)
value MINCHAR (0x80)
value MINIMUM_RESERVED_MANIFEST_RESOURCE_ID (MAKEINTRESOURCE( 1 ))
value MINLONG (0x80000000)
value MINSHORT (0x8000)
value MIN_ACL_REVISION (ACL_REVISION2)
value MIN_LOGICALDPIOVERRIDE (-2)
value MIN_PRIORITY (1)
value MIN_UCSCHAR ((0))
value MIXERCONTROL_CONTROLF_DISABLED (0x80000000L)
value MIXERCONTROL_CONTROLF_MULTIPLE (0x00000002L)
value MIXERCONTROL_CONTROLF_UNIFORM (0x00000001L)
value MIXERCONTROL_CONTROLTYPE_BASS ((MIXERCONTROL_CONTROLTYPE_FADER + 2))
value MIXERCONTROL_CONTROLTYPE_BASS_BOOST ((MIXERCONTROL_CONTROLTYPE_BOOLEAN + 0x00002277))
value MIXERCONTROL_CONTROLTYPE_BOOLEAN ((MIXERCONTROL_CT_CLASS_SWITCH | MIXERCONTROL_CT_SC_SWITCH_BOOLEAN | MIXERCONTROL_CT_UNITS_BOOLEAN))
value MIXERCONTROL_CONTROLTYPE_BOOLEANMETER ((MIXERCONTROL_CT_CLASS_METER | MIXERCONTROL_CT_SC_METER_POLLED | MIXERCONTROL_CT_UNITS_BOOLEAN))
value MIXERCONTROL_CONTROLTYPE_BUTTON ((MIXERCONTROL_CT_CLASS_SWITCH | MIXERCONTROL_CT_SC_SWITCH_BUTTON | MIXERCONTROL_CT_UNITS_BOOLEAN))
value MIXERCONTROL_CONTROLTYPE_CUSTOM ((MIXERCONTROL_CT_CLASS_CUSTOM | MIXERCONTROL_CT_UNITS_CUSTOM))
value MIXERCONTROL_CONTROLTYPE_DECIBELS ((MIXERCONTROL_CT_CLASS_NUMBER | MIXERCONTROL_CT_UNITS_DECIBELS))
value MIXERCONTROL_CONTROLTYPE_EQUALIZER ((MIXERCONTROL_CONTROLTYPE_FADER + 4))
value MIXERCONTROL_CONTROLTYPE_FADER ((MIXERCONTROL_CT_CLASS_FADER | MIXERCONTROL_CT_UNITS_UNSIGNED))
value MIXERCONTROL_CONTROLTYPE_LOUDNESS ((MIXERCONTROL_CONTROLTYPE_BOOLEAN + 4))
value MIXERCONTROL_CONTROLTYPE_MICROTIME ((MIXERCONTROL_CT_CLASS_TIME | MIXERCONTROL_CT_SC_TIME_MICROSECS | MIXERCONTROL_CT_UNITS_UNSIGNED))
value MIXERCONTROL_CONTROLTYPE_MILLITIME ((MIXERCONTROL_CT_CLASS_TIME | MIXERCONTROL_CT_SC_TIME_MILLISECS | MIXERCONTROL_CT_UNITS_UNSIGNED))
value MIXERCONTROL_CONTROLTYPE_MIXER ((MIXERCONTROL_CONTROLTYPE_MULTIPLESELECT + 1))
value MIXERCONTROL_CONTROLTYPE_MONO ((MIXERCONTROL_CONTROLTYPE_BOOLEAN + 3))
value MIXERCONTROL_CONTROLTYPE_MULTIPLESELECT ((MIXERCONTROL_CT_CLASS_LIST | MIXERCONTROL_CT_SC_LIST_MULTIPLE | MIXERCONTROL_CT_UNITS_BOOLEAN))
value MIXERCONTROL_CONTROLTYPE_MUTE ((MIXERCONTROL_CONTROLTYPE_BOOLEAN + 2))
value MIXERCONTROL_CONTROLTYPE_MUX ((MIXERCONTROL_CONTROLTYPE_SINGLESELECT + 1))
value MIXERCONTROL_CONTROLTYPE_ONOFF ((MIXERCONTROL_CONTROLTYPE_BOOLEAN + 1))
value MIXERCONTROL_CONTROLTYPE_PAN ((MIXERCONTROL_CONTROLTYPE_SLIDER + 1))
value MIXERCONTROL_CONTROLTYPE_PEAKMETER ((MIXERCONTROL_CONTROLTYPE_SIGNEDMETER + 1))
value MIXERCONTROL_CONTROLTYPE_PERCENT ((MIXERCONTROL_CT_CLASS_NUMBER | MIXERCONTROL_CT_UNITS_PERCENT))
value MIXERCONTROL_CONTROLTYPE_QSOUNDPAN ((MIXERCONTROL_CONTROLTYPE_SLIDER + 2))
value MIXERCONTROL_CONTROLTYPE_SIGNED ((MIXERCONTROL_CT_CLASS_NUMBER | MIXERCONTROL_CT_UNITS_SIGNED))
value MIXERCONTROL_CONTROLTYPE_SIGNEDMETER ((MIXERCONTROL_CT_CLASS_METER | MIXERCONTROL_CT_SC_METER_POLLED | MIXERCONTROL_CT_UNITS_SIGNED))
value MIXERCONTROL_CONTROLTYPE_SINGLESELECT ((MIXERCONTROL_CT_CLASS_LIST | MIXERCONTROL_CT_SC_LIST_SINGLE | MIXERCONTROL_CT_UNITS_BOOLEAN))
value MIXERCONTROL_CONTROLTYPE_SLIDER ((MIXERCONTROL_CT_CLASS_SLIDER | MIXERCONTROL_CT_UNITS_SIGNED))
value MIXERCONTROL_CONTROLTYPE_STEREOENH ((MIXERCONTROL_CONTROLTYPE_BOOLEAN + 5))
value MIXERCONTROL_CONTROLTYPE_TREBLE ((MIXERCONTROL_CONTROLTYPE_FADER + 3))
value MIXERCONTROL_CONTROLTYPE_UNSIGNED ((MIXERCONTROL_CT_CLASS_NUMBER | MIXERCONTROL_CT_UNITS_UNSIGNED))
value MIXERCONTROL_CONTROLTYPE_UNSIGNEDMETER ((MIXERCONTROL_CT_CLASS_METER | MIXERCONTROL_CT_SC_METER_POLLED | MIXERCONTROL_CT_UNITS_UNSIGNED))
value MIXERCONTROL_CONTROLTYPE_VOLUME ((MIXERCONTROL_CONTROLTYPE_FADER + 1))
value MIXERCONTROL_CT_CLASS_CUSTOM (0x00000000L)
value MIXERCONTROL_CT_CLASS_FADER (0x50000000L)
value MIXERCONTROL_CT_CLASS_LIST (0x70000000L)
value MIXERCONTROL_CT_CLASS_MASK (0xF0000000L)
value MIXERCONTROL_CT_CLASS_METER (0x10000000L)
value MIXERCONTROL_CT_CLASS_NUMBER (0x30000000L)
value MIXERCONTROL_CT_CLASS_SLIDER (0x40000000L)
value MIXERCONTROL_CT_CLASS_SWITCH (0x20000000L)
value MIXERCONTROL_CT_CLASS_TIME (0x60000000L)
value MIXERCONTROL_CT_SC_LIST_MULTIPLE (0x01000000L)
value MIXERCONTROL_CT_SC_LIST_SINGLE (0x00000000L)
value MIXERCONTROL_CT_SC_METER_POLLED (0x00000000L)
value MIXERCONTROL_CT_SC_SWITCH_BOOLEAN (0x00000000L)
value MIXERCONTROL_CT_SC_SWITCH_BUTTON (0x01000000L)
value MIXERCONTROL_CT_SC_TIME_MICROSECS (0x00000000L)
value MIXERCONTROL_CT_SC_TIME_MILLISECS (0x01000000L)
value MIXERCONTROL_CT_SUBCLASS_MASK (0x0F000000L)
value MIXERCONTROL_CT_UNITS_BOOLEAN (0x00010000L)
value MIXERCONTROL_CT_UNITS_CUSTOM (0x00000000L)
value MIXERCONTROL_CT_UNITS_DECIBELS (0x00040000L)
value MIXERCONTROL_CT_UNITS_MASK (0x00FF0000L)
value MIXERCONTROL_CT_UNITS_PERCENT (0x00050000L)
value MIXERCONTROL_CT_UNITS_SIGNED (0x00020000L)
value MIXERCONTROL_CT_UNITS_UNSIGNED (0x00030000L)
value MIXERLINE_COMPONENTTYPE_DST_DIGITAL ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 1))
value MIXERLINE_COMPONENTTYPE_DST_FIRST (0x00000000L)
value MIXERLINE_COMPONENTTYPE_DST_HEADPHONES ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 5))
value MIXERLINE_COMPONENTTYPE_DST_LAST ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 8))
value MIXERLINE_COMPONENTTYPE_DST_LINE ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 2))
value MIXERLINE_COMPONENTTYPE_DST_MONITOR ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 3))
value MIXERLINE_COMPONENTTYPE_DST_SPEAKERS ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 4))
value MIXERLINE_COMPONENTTYPE_DST_TELEPHONE ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 6))
value MIXERLINE_COMPONENTTYPE_DST_UNDEFINED ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 0))
value MIXERLINE_COMPONENTTYPE_DST_VOICEIN ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 8))
value MIXERLINE_COMPONENTTYPE_DST_WAVEIN ((MIXERLINE_COMPONENTTYPE_DST_FIRST + 7))
value MIXERLINE_COMPONENTTYPE_SRC_ANALOG ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 10))
value MIXERLINE_COMPONENTTYPE_SRC_AUXILIARY ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 9))
value MIXERLINE_COMPONENTTYPE_SRC_COMPACTDISC ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 5))
value MIXERLINE_COMPONENTTYPE_SRC_DIGITAL ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 1))
value MIXERLINE_COMPONENTTYPE_SRC_FIRST (0x00001000L)
value MIXERLINE_COMPONENTTYPE_SRC_LAST ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 10))
value MIXERLINE_COMPONENTTYPE_SRC_LINE ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 2))
value MIXERLINE_COMPONENTTYPE_SRC_MICROPHONE ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 3))
value MIXERLINE_COMPONENTTYPE_SRC_PCSPEAKER ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 7))
value MIXERLINE_COMPONENTTYPE_SRC_SYNTHESIZER ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 4))
value MIXERLINE_COMPONENTTYPE_SRC_TELEPHONE ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 6))
value MIXERLINE_COMPONENTTYPE_SRC_UNDEFINED ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 0))
value MIXERLINE_COMPONENTTYPE_SRC_WAVEOUT ((MIXERLINE_COMPONENTTYPE_SRC_FIRST + 8))
value MIXERLINE_LINEF_ACTIVE (0x00000001L)
value MIXERLINE_LINEF_DISCONNECTED (0x00008000L)
value MIXERLINE_LINEF_SOURCE (0x80000000L)
value MIXERLINE_TARGETTYPE_AUX (5)
value MIXERLINE_TARGETTYPE_MIDIIN (4)
value MIXERLINE_TARGETTYPE_MIDIOUT (3)
value MIXERLINE_TARGETTYPE_UNDEFINED (0)
value MIXERLINE_TARGETTYPE_WAVEIN (2)
value MIXERLINE_TARGETTYPE_WAVEOUT (1)
value MIXERR_BASE (1024)
value MIXERR_INVALCONTROL ((MIXERR_BASE + 1))
value MIXERR_INVALLINE ((MIXERR_BASE + 0))
value MIXERR_INVALVALUE ((MIXERR_BASE + 2))
value MIXERR_LASTERROR ((MIXERR_BASE + 2))
value MIXER_GETCONTROLDETAILSF_LISTTEXT (0x00000001L)
value MIXER_GETCONTROLDETAILSF_QUERYMASK (0x0000000FL)
value MIXER_GETCONTROLDETAILSF_VALUE (0x00000000L)
value MIXER_GETLINECONTROLSF_ALL (0x00000000L)
value MIXER_GETLINECONTROLSF_ONEBYID (0x00000001L)
value MIXER_GETLINECONTROLSF_ONEBYTYPE (0x00000002L)
value MIXER_GETLINECONTROLSF_QUERYMASK (0x0000000FL)
value MIXER_GETLINEINFOF_COMPONENTTYPE (0x00000003L)
value MIXER_GETLINEINFOF_DESTINATION (0x00000000L)
value MIXER_GETLINEINFOF_LINEID (0x00000002L)
value MIXER_GETLINEINFOF_QUERYMASK (0x0000000FL)
value MIXER_GETLINEINFOF_SOURCE (0x00000001L)
value MIXER_GETLINEINFOF_TARGETTYPE (0x00000004L)
value MIXER_LONG_NAME_CHARS (64)
value MIXER_OBJECTF_AUX (0x50000000L)
value MIXER_OBJECTF_HANDLE (0x80000000L)
value MIXER_OBJECTF_HMIDIIN ((MIXER_OBJECTF_HANDLE|MIXER_OBJECTF_MIDIIN))
value MIXER_OBJECTF_HMIDIOUT ((MIXER_OBJECTF_HANDLE|MIXER_OBJECTF_MIDIOUT))
value MIXER_OBJECTF_HMIXER ((MIXER_OBJECTF_HANDLE|MIXER_OBJECTF_MIXER))
value MIXER_OBJECTF_HWAVEIN ((MIXER_OBJECTF_HANDLE|MIXER_OBJECTF_WAVEIN))
value MIXER_OBJECTF_HWAVEOUT ((MIXER_OBJECTF_HANDLE|MIXER_OBJECTF_WAVEOUT))
value MIXER_OBJECTF_MIDIIN (0x40000000L)
value MIXER_OBJECTF_MIDIOUT (0x30000000L)
value MIXER_OBJECTF_MIXER (0x00000000L)
value MIXER_OBJECTF_WAVEIN (0x20000000L)
value MIXER_OBJECTF_WAVEOUT (0x10000000L)
value MIXER_SETCONTROLDETAILSF_CUSTOM (0x00000001L)
value MIXER_SETCONTROLDETAILSF_QUERYMASK (0x0000000FL)
value MIXER_SETCONTROLDETAILSF_VALUE (0x00000000L)
value MIXER_SHORT_NAME_CHARS (16)
value MKF_AVAILABLE (0x00000002)
value MKF_CONFIRMHOTKEY (0x00000008)
value MKF_HOTKEYACTIVE (0x00000004)
value MKF_HOTKEYSOUND (0x00000010)
value MKF_INDICATOR (0x00000020)
value MKF_LEFTBUTTONDOWN (0x01000000)
value MKF_LEFTBUTTONSEL (0x10000000)
value MKF_MODIFIERS (0x00000040)
value MKF_MOUSEKEYSON (0x00000001)
value MKF_MOUSEMODE (0x80000000)
value MKF_REPLACENUMBERS (0x00000080)
value MKF_RIGHTBUTTONDOWN (0x02000000)
value MKF_RIGHTBUTTONSEL (0x20000000)
value MKSYS_URLMONIKER (6)
value MK_ALT (( 0x20 ))
value MK_CONTROL (0x0008)
value MK_E_CANTOPENFILE (_HRESULT_TYPEDEF_(0x800401EAL))
value MK_E_CONNECTMANUALLY (_HRESULT_TYPEDEF_(0x800401E0L))
value MK_E_ENUMERATION_FAILED (_HRESULT_TYPEDEF_(0x800401EFL))
value MK_E_EXCEEDEDDEADLINE (_HRESULT_TYPEDEF_(0x800401E1L))
value MK_E_FIRST (0x800401E0L)
value MK_E_INTERMEDIATEINTERFACENOTSUPPORTED (_HRESULT_TYPEDEF_(0x800401E7L))
value MK_E_INVALIDEXTENSION (_HRESULT_TYPEDEF_(0x800401E6L))
value MK_E_LAST (0x800401EFL)
value MK_E_MUSTBOTHERUSER (_HRESULT_TYPEDEF_(0x800401EBL))
value MK_E_NEEDGENERIC (_HRESULT_TYPEDEF_(0x800401E2L))
value MK_E_NOINVERSE (_HRESULT_TYPEDEF_(0x800401ECL))
value MK_E_NOOBJECT (_HRESULT_TYPEDEF_(0x800401E5L))
value MK_E_NOPREFIX (_HRESULT_TYPEDEF_(0x800401EEL))
value MK_E_NOSTORAGE (_HRESULT_TYPEDEF_(0x800401EDL))
value MK_E_NOTBINDABLE (_HRESULT_TYPEDEF_(0x800401E8L))
value MK_E_NOTBOUND (_HRESULT_TYPEDEF_(0x800401E9L))
value MK_E_NO_NORMALIZED (_HRESULT_TYPEDEF_(0x80080007L))
value MK_E_SYNTAX (_HRESULT_TYPEDEF_(0x800401E4L))
value MK_E_UNAVAILABLE (_HRESULT_TYPEDEF_(0x800401E3L))
value MK_LBUTTON (0x0001)
value MK_MBUTTON (0x0010)
value MK_RBUTTON (0x0002)
value MK_SHIFT (0x0004)
value MK_S_ASYNCHRONOUS (_HRESULT_TYPEDEF_(0x000401E8L))
value MK_S_FIRST (0x000401E0L)
value MK_S_HIM (_HRESULT_TYPEDEF_(0x000401E5L))
value MK_S_LAST (0x000401EFL)
value MK_S_ME (_HRESULT_TYPEDEF_(0x000401E4L))
value MK_S_MONIKERALREADYREGISTERED (_HRESULT_TYPEDEF_(0x000401E7L))
value MK_S_REDUCED_TO_SELF (_HRESULT_TYPEDEF_(0x000401E2L))
value MK_S_US (_HRESULT_TYPEDEF_(0x000401E6L))
value MMIOERR_ACCESSDENIED ((MMIOERR_BASE + 12))
value MMIOERR_BASE (256)
value MMIOERR_CANNOTCLOSE ((MMIOERR_BASE + 4))
value MMIOERR_CANNOTEXPAND ((MMIOERR_BASE + 8))
value MMIOERR_CANNOTOPEN ((MMIOERR_BASE + 3))
value MMIOERR_CANNOTREAD ((MMIOERR_BASE + 5))
value MMIOERR_CANNOTSEEK ((MMIOERR_BASE + 7))
value MMIOERR_CANNOTWRITE ((MMIOERR_BASE + 6))
value MMIOERR_CHUNKNOTFOUND ((MMIOERR_BASE + 9))
value MMIOERR_FILENOTFOUND ((MMIOERR_BASE + 1))
value MMIOERR_INVALIDFILE ((MMIOERR_BASE + 16))
value MMIOERR_NETWORKERROR ((MMIOERR_BASE + 14))
value MMIOERR_OUTOFMEMORY ((MMIOERR_BASE + 2))
value MMIOERR_PATHNOTFOUND ((MMIOERR_BASE + 11))
value MMIOERR_SHARINGVIOLATION ((MMIOERR_BASE + 13))
value MMIOERR_TOOMANYOPENFILES ((MMIOERR_BASE + 15))
value MMIOERR_UNBUFFERED ((MMIOERR_BASE + 10))
value MMIOM_CLOSE (4)
value MMIOM_OPEN (3)
value MMIOM_READ (MMIO_READ)
value MMIOM_RENAME (6)
value MMIOM_SEEK (2)
value MMIOM_USER (0x8000)
value MMIOM_WRITE (MMIO_WRITE)
value MMIOM_WRITEFLUSH (5)
value MMIO_ALLOCBUF (0x00010000)
value MMIO_COMPAT (0x00000000)
value MMIO_CREATE (0x00001000)
value MMIO_CREATELIST (0x0040)
value MMIO_CREATERIFF (0x0020)
value MMIO_DEFAULTBUFFER (8192)
value MMIO_DELETE (0x00000200)
value MMIO_DENYNONE (0x00000040)
value MMIO_DENYREAD (0x00000030)
value MMIO_DENYWRITE (0x00000020)
value MMIO_DIRTY (0x10000000)
value MMIO_EMPTYBUF (0x0010)
value MMIO_EXCLUSIVE (0x00000010)
value MMIO_EXIST (0x00004000)
value MMIO_FHOPEN (0x0010)
value MMIO_FINDCHUNK (0x0010)
value MMIO_FINDLIST (0x0040)
value MMIO_FINDPROC (0x00040000)
value MMIO_FINDRIFF (0x0020)
value MMIO_GETTEMP (0x00020000)
value MMIO_GLOBALPROC (0x10000000)
value MMIO_INSTALLPROC (0x00010000)
value MMIO_PARSE (0x00000100)
value MMIO_READ (0x00000000)
value MMIO_READWRITE (0x00000002)
value MMIO_REMOVEPROC (0x00020000)
value MMIO_RWMODE (0x00000003)
value MMIO_SHAREMODE (0x00000070)
value MMIO_TOUPPER (0x0010)
value MMIO_UNICODEPROC (0x01000000)
value MMIO_WRITE (0x00000001)
value MMSYSERR_ALLOCATED ((MMSYSERR_BASE + 4))
value MMSYSERR_BADDB ((MMSYSERR_BASE + 14))
value MMSYSERR_BADDEVICEID ((MMSYSERR_BASE + 2))
value MMSYSERR_BADERRNUM ((MMSYSERR_BASE + 9))
value MMSYSERR_BASE (0)
value MMSYSERR_DELETEERROR ((MMSYSERR_BASE + 18))
value MMSYSERR_ERROR ((MMSYSERR_BASE + 1))
value MMSYSERR_HANDLEBUSY ((MMSYSERR_BASE + 12))
value MMSYSERR_INVALFLAG ((MMSYSERR_BASE + 10))
value MMSYSERR_INVALHANDLE ((MMSYSERR_BASE + 5))
value MMSYSERR_INVALIDALIAS ((MMSYSERR_BASE + 13))
value MMSYSERR_INVALPARAM ((MMSYSERR_BASE + 11))
value MMSYSERR_KEYNOTFOUND ((MMSYSERR_BASE + 15))
value MMSYSERR_LASTERROR ((MMSYSERR_BASE + 21))
value MMSYSERR_MOREDATA ((MMSYSERR_BASE + 21))
value MMSYSERR_NODRIVER ((MMSYSERR_BASE + 6))
value MMSYSERR_NODRIVERCB ((MMSYSERR_BASE + 20))
value MMSYSERR_NOERROR (0)
value MMSYSERR_NOMEM ((MMSYSERR_BASE + 7))
value MMSYSERR_NOTENABLED ((MMSYSERR_BASE + 3))
value MMSYSERR_NOTSUPPORTED ((MMSYSERR_BASE + 8))
value MMSYSERR_READERROR ((MMSYSERR_BASE + 16))
value MMSYSERR_VALNOTFOUND ((MMSYSERR_BASE + 19))
value MMSYSERR_WRITEERROR ((MMSYSERR_BASE + 17))
value MM_ANISOTROPIC (8)
value MM_DRVM_CLOSE (0x3D1)
value MM_DRVM_DATA (0x3D2)
value MM_DRVM_ERROR (0x3D3)
value MM_DRVM_OPEN (0x3D0)
value MM_HIENGLISH (5)
value MM_HIMETRIC (3)
value MM_ISOTROPIC (7)
value MM_LOENGLISH (4)
value MM_LOMETRIC (2)
value MM_MAX (MM_ANISOTROPIC)
value MM_MAX_AXES_NAMELEN (16)
value MM_MAX_FIXEDSCALE (MM_TWIPS)
value MM_MAX_NUMAXES (16)
value MM_MCINOTIFY (0x3B9)
value MM_MCISIGNAL (0x3CB)
value MM_MIM_CLOSE (0x3C2)
value MM_MIM_DATA (0x3C3)
value MM_MIM_ERROR (0x3C5)
value MM_MIM_LONGDATA (0x3C4)
value MM_MIM_LONGERROR (0x3C6)
value MM_MIM_MOREDATA (0x3CC)
value MM_MIM_OPEN (0x3C1)
value MM_MIN (MM_TEXT)
value MM_MIXM_CONTROL_CHANGE (0x3D1)
value MM_MIXM_LINE_CHANGE (0x3D0)
value MM_MOM_CLOSE (0x3C8)
value MM_MOM_DONE (0x3C9)
value MM_MOM_OPEN (0x3C7)
value MM_MOM_POSITIONCB (0x3CA)
value MM_STREAM_CLOSE (0x3D5)
value MM_STREAM_DONE (0x3D6)
value MM_STREAM_ERROR (0x3D7)
value MM_STREAM_OPEN (0x3D4)
value MM_TEXT (1)
value MM_TWIPS (6)
value MM_WIM_CLOSE (0x3BF)
value MM_WIM_DATA (0x3C0)
value MM_WIM_OPEN (0x3BE)
value MM_WOM_CLOSE (0x3BC)
value MM_WOM_DONE (0x3BD)
value MM_WOM_OPEN (0x3BB)
value MNC_CLOSE (1)
value MNC_EXECUTE (2)
value MNC_IGNORE (0)
value MNC_SELECT (3)
value MND_CONTINUE (0)
value MND_ENDMENU (1)
value MNGOF_BOTTOMGAP (0x00000002)
value MNGOF_TOPGAP (0x00000001)
value MNGO_NOERROR (0x00000001)
value MNGO_NOINTERFACE (0x00000000)
value MNS_AUTODISMISS (0x10000000)
value MNS_CHECKORBMP (0x04000000)
value MNS_DRAGDROP (0x20000000)
value MNS_MODELESS (0x40000000)
value MNS_NOCHECK (0x80000000)
value MNS_NOTIFYBYPOS (0x08000000)
value MN_GETHMENU (0x01E1)
value MOD_ALT (0x0001)
value MOD_CONTROL (0x0002)
value MOD_FMSYNTH (4)
value MOD_IGNORE_ALL_MODIFIER (0x0400)
value MOD_LEFT (0x8000)
value MOD_MAPPER (5)
value MOD_MIDIPORT (1)
value MOD_NOREPEAT (0x4000)
value MOD_ON_KEYUP (0x0800)
value MOD_RIGHT (0x4000)
value MOD_SHIFT (0x0004)
value MOD_SQSYNTH (3)
value MOD_SWSYNTH (7)
value MOD_SYNTH (2)
value MOD_WAVETABLE (6)
value MOD_WIN (0x0008)
value MOM_CLOSE (MM_MOM_CLOSE)
value MOM_DONE (MM_MOM_DONE)
value MOM_OPEN (MM_MOM_OPEN)
value MOM_POSITIONCB (MM_MOM_POSITIONCB)
value MONITORINFOF_PRIMARY (0x00000001)
value MONITOR_DEFAULTTONEAREST (0x00000002)
value MONITOR_DEFAULTTONULL (0x00000000)
value MONITOR_DEFAULTTOPRIMARY (0x00000001)
value MONO_FONT (8)
value MOUSEEVENTF_ABSOLUTE (0x8000)
value MOUSEEVENTF_HWHEEL (0x01000)
value MOUSEEVENTF_LEFTDOWN (0x0002)
value MOUSEEVENTF_LEFTUP (0x0004)
value MOUSEEVENTF_MIDDLEDOWN (0x0020)
value MOUSEEVENTF_MIDDLEUP (0x0040)
value MOUSEEVENTF_MOVE (0x0001)
value MOUSEEVENTF_MOVE_NOCOALESCE (0x2000)
value MOUSEEVENTF_RIGHTDOWN (0x0008)
value MOUSEEVENTF_RIGHTUP (0x0010)
value MOUSEEVENTF_VIRTUALDESK (0x4000)
value MOUSEEVENTF_WHEEL (0x0800)
value MOUSEEVENTF_XDOWN (0x0080)
value MOUSEEVENTF_XUP (0x0100)
value MOUSETRAILS (39)
value MOUSEWHEEL_ROUTING_FOCUS (0)
value MOUSEWHEEL_ROUTING_HYBRID (1)
value MOUSEWHEEL_ROUTING_MOUSE_POS (2)
value MOUSE_ATTRIBUTES_CHANGED (0x04)
value MOUSE_EVENT (0x0002)
value MOUSE_HWHEELED (0x0008)
value MOUSE_MOVED (0x0001)
value MOUSE_MOVE_ABSOLUTE (1)
value MOUSE_MOVE_NOCOALESCE (0x08)
value MOUSE_MOVE_RELATIVE (0)
value MOUSE_VIRTUAL_DESKTOP (0x02)
value MOUSE_WHEELED (0x0004)
value MOVEFILE_COPY_ALLOWED (0x00000002)
value MOVEFILE_CREATE_HARDLINK (0x00000010)
value MOVEFILE_DELAY_UNTIL_REBOOT (0x00000004)
value MOVEFILE_FAIL_IF_NOT_TRACKABLE (0x00000020)
value MOVEFILE_REPLACE_EXISTING (0x00000001)
value MOVEFILE_WRITE_THROUGH (0x00000008)
value MSDTC_E_DUPLICATE_RESOURCE (_HRESULT_TYPEDEF_(0x80110701L))
value MSGFLTINFO_ALLOWED_HIGHER ((3))
value MSGFLTINFO_ALREADYALLOWED_FORWND ((1))
value MSGFLTINFO_ALREADYDISALLOWED_FORWND ((2))
value MSGFLTINFO_NONE ((0))
value MSGFLT_ADD (1)
value MSGFLT_ALLOW ((1))
value MSGFLT_DISALLOW ((2))
value MSGFLT_REMOVE (2)
value MSGFLT_RESET ((0))
value MSGF_DDEMGR (0x8001)
value MSGF_DIALOGBOX (0)
value MSGF_MAX (8)
value MSGF_MENU (2)
value MSGF_MESSAGEBOX (1)
value MSGF_NEXTWINDOW (6)
value MSGF_SCROLLBAR (5)
value MSGF_USER (4096)
value MSG_BCAST (0x0400)
value MSG_CTRUNC (0x0200)
value MSG_DONTROUTE (0x4)
value MSG_ERRQUEUE (0x1000)
value MSG_INTERRUPT (0x10)
value MSG_MAXIOVLEN (16)
value MSG_MCAST (0x0800)
value MSG_OOB (0x1)
value MSG_PARTIAL (0x8000)
value MSG_PEEK (0x2)
value MSG_PUSH_IMMEDIATE (0x20)
value MSG_TRUNC (0x0100)
value MSG_WAITALL (0x8)
value MSSIPOTF_E_BADVERSION (_HRESULT_TYPEDEF_(0x80097015L))
value MSSIPOTF_E_BAD_FIRST_TABLE_PLACEMENT (_HRESULT_TYPEDEF_(0x80097008L))
value MSSIPOTF_E_BAD_MAGICNUMBER (_HRESULT_TYPEDEF_(0x80097004L))
value MSSIPOTF_E_BAD_OFFSET_TABLE (_HRESULT_TYPEDEF_(0x80097005L))
value MSSIPOTF_E_CANTGETOBJECT (_HRESULT_TYPEDEF_(0x80097002L))
value MSSIPOTF_E_CRYPT (_HRESULT_TYPEDEF_(0x80097014L))
value MSSIPOTF_E_DSIG_STRUCTURE (_HRESULT_TYPEDEF_(0x80097016L))
value MSSIPOTF_E_FAILED_HINTS_CHECK (_HRESULT_TYPEDEF_(0x80097011L))
value MSSIPOTF_E_FAILED_POLICY (_HRESULT_TYPEDEF_(0x80097010L))
value MSSIPOTF_E_FILE (_HRESULT_TYPEDEF_(0x80097013L))
value MSSIPOTF_E_FILETOOSMALL (_HRESULT_TYPEDEF_(0x8009700BL))
value MSSIPOTF_E_FILE_CHECKSUM (_HRESULT_TYPEDEF_(0x8009700DL))
value MSSIPOTF_E_NOHEADTABLE (_HRESULT_TYPEDEF_(0x80097003L))
value MSSIPOTF_E_NOT_OPENTYPE (_HRESULT_TYPEDEF_(0x80097012L))
value MSSIPOTF_E_OUTOFMEMRANGE (_HRESULT_TYPEDEF_(0x80097001L))
value MSSIPOTF_E_PCONST_CHECK (_HRESULT_TYPEDEF_(0x80097017L))
value MSSIPOTF_E_STRUCTURE (_HRESULT_TYPEDEF_(0x80097018L))
value MSSIPOTF_E_TABLES_OVERLAP (_HRESULT_TYPEDEF_(0x80097009L))
value MSSIPOTF_E_TABLE_CHECKSUM (_HRESULT_TYPEDEF_(0x8009700CL))
value MSSIPOTF_E_TABLE_LONGWORD (_HRESULT_TYPEDEF_(0x80097007L))
value MSSIPOTF_E_TABLE_PADBYTES (_HRESULT_TYPEDEF_(0x8009700AL))
value MSSIPOTF_E_TABLE_TAGORDER (_HRESULT_TYPEDEF_(0x80097006L))
value MS_CTS_ON (((DWORD)0x0010))
value MS_DEF_DH_SCHANNEL_PROV (MS_DEF_DH_SCHANNEL_PROV_A)
value MS_DEF_DSS_DH_PROV (MS_DEF_DSS_DH_PROV_A)
value MS_DEF_DSS_PROV (MS_DEF_DSS_PROV_A)
value MS_DEF_PROV (MS_DEF_PROV_A)
value MS_DEF_RSA_SCHANNEL_PROV (MS_DEF_RSA_SCHANNEL_PROV_A)
value MS_DEF_RSA_SIG_PROV (MS_DEF_RSA_SIG_PROV_A)
value MS_DSR_ON (((DWORD)0x0020))
value MS_ENHANCED_PROV (MS_ENHANCED_PROV_A)
value MS_ENH_DSS_DH_PROV (MS_ENH_DSS_DH_PROV_A)
value MS_ENH_RSA_AES_PROV (MS_ENH_RSA_AES_PROV_A)
value MS_ENH_RSA_AES_PROV_XP (MS_ENH_RSA_AES_PROV_XP_A)
value MS_PPM_SOFTWARE_ALL (0x1)
value MS_RING_ON (((DWORD)0x0040))
value MS_RLSD_ON (((DWORD)0x0080))
value MS_SCARD_PROV (MS_SCARD_PROV_A)
value MS_STRONG_PROV (MS_STRONG_PROV_A)
value MUI_CALLBACK_ALL_FLAGS (MUI_CALLBACK_FLAG_UPGRADED_INSTALLATION)
value MUI_COMPLEX_SCRIPT_FILTER (0x200)
value MUI_CONSOLE_FILTER (0x100)
value MUI_FILEINFO_VERSION (0x001)
value MUI_FILETYPE_LANGUAGE_NEUTRAL_MAIN (0x002)
value MUI_FILETYPE_LANGUAGE_NEUTRAL_MUI (0x004)
value MUI_FILETYPE_NOT_LANGUAGE_NEUTRAL (0x001)
value MUI_FORMAT_INF_COMPAT (0x0002)
value MUI_FORMAT_REG_COMPAT (0x0001)
value MUI_FULL_LANGUAGE (0x01)
value MUI_IMMUTABLE_LOOKUP (0x0010)
value MUI_LANGUAGE_ID (0x4)
value MUI_LANGUAGE_INSTALLED (0x20)
value MUI_LANGUAGE_LICENSED (0x40)
value MUI_LANGUAGE_NAME (0x8)
value MUI_LANG_NEUTRAL_PE_FILE (0x100)
value MUI_LIP_LANGUAGE (0x04)
value MUI_MACHINE_LANGUAGE_SETTINGS (0x400)
value MUI_MERGE_SYSTEM_FALLBACK (0x10)
value MUI_MERGE_USER_FALLBACK (0x20)
value MUI_NON_LANG_NEUTRAL_FILE (0x200)
value MUI_PARTIAL_LANGUAGE (0x02)
value MUI_QUERY_CHECKSUM (0x002)
value MUI_QUERY_LANGUAGE_NAME (0x004)
value MUI_QUERY_RESOURCE_TYPES (0x008)
value MUI_QUERY_TYPE (0x001)
value MUI_RESET_FILTERS (0x001)
value MUI_SKIP_STRING_CACHE (0x0008)
value MUI_THREAD_LANGUAGES (0x40)
value MUI_UI_FALLBACK (MUI_MERGE_SYSTEM_FALLBACK | MUI_MERGE_USER_FALLBACK)
value MUI_USER_PREFERRED_UI_LANGUAGES (0x10)
value MUI_USE_INSTALLED_LANGUAGES (0x20)
value MUI_USE_SEARCH_ALL_LANGUAGES (0x40)
value MUI_VERIFY_FILE_EXISTS (0x0004)
value MULTIFILEOPENORD (1537)
value MUTANT_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED|SYNCHRONIZE| MUTANT_QUERY_STATE))
value MUTANT_QUERY_STATE (0x0001)
value MUTEX_ALL_ACCESS (MUTANT_ALL_ACCESS)
value MUTEX_MODIFY_STATE (MUTANT_QUERY_STATE)
value MUTZ_ACCEPT_WILDCARD_SCHEME (0x00000080)
value MUTZ_DONT_UNESCAPE (0x00000800)
value MUTZ_DONT_USE_CACHE (0x00001000)
value MUTZ_ENFORCERESTRICTED (0x00000100)
value MUTZ_FORCE_INTRANET_FLAGS (0x00002000)
value MUTZ_IGNORE_ZONE_MAPPINGS (0x00004000)
value MUTZ_ISFILE (0x00000002)
value MUTZ_NOSAVEDFILECHECK (0x00000001)
value MUTZ_REQUIRESAVEDFILECHECK (0x00000400)
value MUTZ_RESERVED (0x00000200)
value MWMO_ALERTABLE (0x0002)
value MWMO_INPUTAVAILABLE (0x0004)
value MWMO_WAITALL (0x0001)
value MWT_IDENTITY (1)
value MWT_LEFTMULTIPLY (2)
value MWT_MAX (MWT_RIGHTMULTIPLY)
value MWT_MIN (MWT_IDENTITY)
value MWT_RIGHTMULTIPLY (3)
value NAME_FLAGS_MASK (0x87)
value NAP_E_CONFLICTING_ID (_HRESULT_TYPEDEF_(0x80270003L))
value NAP_E_ENTITY_DISABLED (_HRESULT_TYPEDEF_(0x8027000EL))
value NAP_E_ID_NOT_FOUND (_HRESULT_TYPEDEF_(0x8027000AL))
value NAP_E_INVALID_PACKET (_HRESULT_TYPEDEF_(0x80270001L))
value NAP_E_MAXSIZE_TOO_SMALL (_HRESULT_TYPEDEF_(0x8027000BL))
value NAP_E_MISMATCHED_ID (_HRESULT_TYPEDEF_(0x80270008L))
value NAP_E_MISSING_SOH (_HRESULT_TYPEDEF_(0x80270002L))
value NAP_E_NETSH_GROUPPOLICY_ERROR (_HRESULT_TYPEDEF_(0x8027000FL))
value NAP_E_NOT_INITIALIZED (_HRESULT_TYPEDEF_(0x80270007L))
value NAP_E_NOT_PENDING (_HRESULT_TYPEDEF_(0x80270009L))
value NAP_E_NOT_REGISTERED (_HRESULT_TYPEDEF_(0x80270006L))
value NAP_E_NO_CACHED_SOH (_HRESULT_TYPEDEF_(0x80270004L))
value NAP_E_SERVICE_NOT_RUNNING (_HRESULT_TYPEDEF_(0x8027000CL))
value NAP_E_SHV_CONFIG_EXISTED (_HRESULT_TYPEDEF_(0x80270011L))
value NAP_E_SHV_CONFIG_NOT_FOUND (_HRESULT_TYPEDEF_(0x80270012L))
value NAP_E_SHV_TIMEOUT (_HRESULT_TYPEDEF_(0x80270013L))
value NAP_E_STILL_BOUND (_HRESULT_TYPEDEF_(0x80270005L))
value NAP_E_TOO_MANY_CALLS (_HRESULT_TYPEDEF_(0x80270010L))
value NAP_S_CERT_ALREADY_PRESENT (_HRESULT_TYPEDEF_(0x0027000DL))
value NCBACTION (0x77)
value NCBADDGRNAME (0x36)
value NCBADDNAME (0x30)
value NCBASTAT (0x33)
value NCBCALL (0x10)
value NCBCANCEL (0x35)
value NCBCHAINSEND (0x17)
value NCBCHAINSENDNA (0x72)
value NCBDELNAME (0x31)
value NCBDGRECV (0x21)
value NCBDGRECVBC (0x23)
value NCBDGSEND (0x20)
value NCBDGSENDBC (0x22)
value NCBENUM (0x37)
value NCBFINDNAME (0x78)
value NCBHANGUP (0x12)
value NCBLANSTALERT (0x73)
value NCBLISTEN (0x11)
value NCBNAMSZ (16)
value NCBRECV (0x15)
value NCBRECVANY (0x16)
value NCBRESET (0x32)
value NCBSEND (0x14)
value NCBSENDNA (0x71)
value NCBSSTAT (0x34)
value NCBTRACE (0x79)
value NCBUNLINK (0x70)
value NCM_DISPLAYERRORTIP ((WM_USER+4))
value NCM_GETADDRESS ((WM_USER+1))
value NCM_GETALLOWTYPE ((WM_USER+3))
value NCM_SETALLOWTYPE ((WM_USER+2))
value NCRYPTBUFFER_ATTESTATIONSTATEMENT_BLOB (51)
value NCRYPTBUFFER_ATTESTATION_CLAIM_CHALLENGE_REQUIRED (53)
value NCRYPTBUFFER_ATTESTATION_CLAIM_TYPE (52)
value NCRYPTBUFFER_CERT_BLOB (47)
value NCRYPTBUFFER_CLAIM_IDBINDING_NONCE (48)
value NCRYPTBUFFER_CLAIM_KEYATTESTATION_NONCE (49)
value NCRYPTBUFFER_DATA (1)
value NCRYPTBUFFER_ECC_CURVE_NAME (60)
value NCRYPTBUFFER_ECC_PARAMETERS (61)
value NCRYPTBUFFER_EMPTY (0)
value NCRYPTBUFFER_KEY_PROPERTY_FLAGS (50)
value NCRYPTBUFFER_PKCS_ALG_ID (43)
value NCRYPTBUFFER_PKCS_ALG_OID (41)
value NCRYPTBUFFER_PKCS_ALG_PARAM (42)
value NCRYPTBUFFER_PKCS_ATTRS (44)
value NCRYPTBUFFER_PKCS_KEY_NAME (45)
value NCRYPTBUFFER_PKCS_OID (40)
value NCRYPTBUFFER_PKCS_SECRET (46)
value NCRYPTBUFFER_PROTECTION_DESCRIPTOR_STRING (3)
value NCRYPTBUFFER_PROTECTION_FLAGS (4)
value NCRYPTBUFFER_SSL_CLEAR_KEY (23)
value NCRYPTBUFFER_SSL_CLIENT_RANDOM (20)
value NCRYPTBUFFER_SSL_HIGHEST_VERSION (22)
value NCRYPTBUFFER_SSL_KEY_ARG_DATA (24)
value NCRYPTBUFFER_SSL_SERVER_RANDOM (21)
value NCRYPTBUFFER_SSL_SESSION_HASH (25)
value NCRYPTBUFFER_TPM_PLATFORM_CLAIM_NONCE (81)
value NCRYPTBUFFER_TPM_PLATFORM_CLAIM_PCR_MASK (80)
value NCRYPTBUFFER_TPM_PLATFORM_CLAIM_STATIC_CREATE (82)
value NCRYPTBUFFER_TPM_SEAL_NO_DA_PROTECTION (73)
value NCRYPTBUFFER_TPM_SEAL_PASSWORD (70)
value NCRYPTBUFFER_TPM_SEAL_POLICYINFO (71)
value NCRYPTBUFFER_TPM_SEAL_TICKET (72)
value NCRYPTBUFFER_VERSION (0)
value NCRYPTBUFFER_VSM_KEY_ATTESTATION_CLAIM_RESTRICTIONS (54)
value NCRYPT_AES_ALGORITHM (BCRYPT_AES_ALGORITHM)
value NCRYPT_AES_ALGORITHM_GROUP (NCRYPT_AES_ALGORITHM)
value NCRYPT_ALLOW_ALL_USAGES (0x00ffffff)
value NCRYPT_ALLOW_ARCHIVING_FLAG (0x00000004)
value NCRYPT_ALLOW_DECRYPT_FLAG (0x00000001)
value NCRYPT_ALLOW_EXPORT_FLAG (0x00000001)
value NCRYPT_ALLOW_KEY_AGREEMENT_FLAG (0x00000004)
value NCRYPT_ALLOW_KEY_IMPORT_FLAG (0x00000008)
value NCRYPT_ALLOW_PLAINTEXT_ARCHIVING_FLAG (0x00000008)
value NCRYPT_ALLOW_PLAINTEXT_EXPORT_FLAG (0x00000002)
value NCRYPT_ALLOW_SIGNING_FLAG (0x00000002)
value NCRYPT_ALLOW_SILENT_KEY_ACCESS (0x00000001)
value NCRYPT_ALTERNATE_KEY_STORAGE_LOCATION_PROPERTY (NCRYPT_PCP_ALTERNATE_KEY_STORAGE_LOCATION_PROPERTY)
value NCRYPT_ASYMMETRIC_ENCRYPTION_INTERFACE (BCRYPT_ASYMMETRIC_ENCRYPTION_INTERFACE)
value NCRYPT_ASYMMETRIC_ENCRYPTION_OPERATION (BCRYPT_ASYMMETRIC_ENCRYPTION_OPERATION)
value NCRYPT_ATTESTATION_FLAG (0x00000020)
value NCRYPT_AUTHORITY_KEY_FLAG (0x00000100)
value NCRYPT_CAPI_KDF_ALGORITHM (BCRYPT_CAPI_KDF_ALGORITHM)
value NCRYPT_CHANGEPASSWORD_PROPERTY (NCRYPT_PCP_CHANGEPASSWORD_PROPERTY)
value NCRYPT_CIPHER_BLOCK_PADDING_FLAG (0x00000001)
value NCRYPT_CIPHER_INTERFACE (BCRYPT_CIPHER_INTERFACE)
value NCRYPT_CIPHER_KEY_BLOB_MAGIC (0x52485043)
value NCRYPT_CIPHER_NO_PADDING_FLAG (0x00000000)
value NCRYPT_CIPHER_OPERATION (BCRYPT_CIPHER_OPERATION)
value NCRYPT_CIPHER_OTHER_PADDING_FLAG (0x00000002)
value NCRYPT_CLAIM_AUTHORITY_AND_SUBJECT (0x00000003)
value NCRYPT_CLAIM_AUTHORITY_ONLY (0x00000001)
value NCRYPT_CLAIM_PLATFORM (0x00010000)
value NCRYPT_CLAIM_SUBJECT_ONLY (0x00000002)
value NCRYPT_CLAIM_UNKNOWN (0x00001000)
value NCRYPT_CLAIM_VSM_KEY_ATTESTATION_STATEMENT (0x00000004)
value NCRYPT_CLAIM_WEB_AUTH_SUBJECT_ONLY (0x00000102)
value NCRYPT_DESX_ALGORITHM (BCRYPT_DESX_ALGORITHM)
value NCRYPT_DES_ALGORITHM (BCRYPT_DES_ALGORITHM)
value NCRYPT_DH_ALGORITHM (BCRYPT_DH_ALGORITHM)
value NCRYPT_DH_ALGORITHM_GROUP (NCRYPT_DH_ALGORITHM)
value NCRYPT_DH_PARAMETERS_PROPERTY (BCRYPT_DH_PARAMETERS)
value NCRYPT_DO_NOT_FINALIZE_FLAG (0x00000400)
value NCRYPT_DSA_ALGORITHM (BCRYPT_DSA_ALGORITHM)
value NCRYPT_DSA_ALGORITHM_GROUP (NCRYPT_DSA_ALGORITHM)
value NCRYPT_ECC_CURVE_NAME_LIST_PROPERTY (BCRYPT_ECC_CURVE_NAME_LIST)
value NCRYPT_ECC_CURVE_NAME_PROPERTY (BCRYPT_ECC_CURVE_NAME)
value NCRYPT_ECC_PARAMETERS_PROPERTY (BCRYPT_ECC_PARAMETERS)
value NCRYPT_ECDH_ALGORITHM (BCRYPT_ECDH_ALGORITHM)
value NCRYPT_ECDSA_ALGORITHM (BCRYPT_ECDSA_ALGORITHM)
value NCRYPT_EXPORTED_ISOLATED_KEY_HEADER_CURRENT_VERSION (NCRYPT_EXPORTED_ISOLATED_KEY_HEADER_V0)
value NCRYPT_EXPORT_LEGACY_FLAG (0x00000800)
value NCRYPT_EXTENDED_ERRORS_FLAG (0x10000000)
value NCRYPT_HASH_INTERFACE (BCRYPT_HASH_INTERFACE)
value NCRYPT_HASH_OPERATION (BCRYPT_HASH_OPERATION)
value NCRYPT_IGNORE_DEVICE_STATE_FLAG (0x00001000)
value NCRYPT_IMPL_HARDWARE_FLAG (0x00000001)
value NCRYPT_IMPL_HARDWARE_RNG_FLAG (0x00000010)
value NCRYPT_IMPL_REMOVABLE_FLAG (0x00000008)
value NCRYPT_IMPL_SOFTWARE_FLAG (0x00000002)
value NCRYPT_IMPL_VIRTUAL_ISOLATION_FLAG (0x00000020)
value NCRYPT_INITIALIZATION_VECTOR (BCRYPT_INITIALIZATION_VECTOR)
value NCRYPT_ISOLATED_KEY_ATTESTED_ATTRIBUTES_CURRENT_VERSION (NCRYPT_ISOLATED_KEY_ATTESTED_ATTRIBUTES_V0)
value NCRYPT_ISOLATED_KEY_FLAG_CREATED_IN_ISOLATION (0x00000001)
value NCRYPT_ISOLATED_KEY_FLAG_IMPORT_ONLY (0x00000002)
value NCRYPT_KDF_KEY_BLOB_MAGIC (0x3146444B)
value NCRYPT_KEY_ACCESS_POLICY_VERSION (1)
value NCRYPT_KEY_ATTEST_MAGIC (0x4450414b)
value NCRYPT_KEY_DERIVATION_INTERFACE (BCRYPT_KEY_DERIVATION_INTERFACE)
value NCRYPT_KEY_DERIVATION_OPERATION (BCRYPT_KEY_DERIVATION_OPERATION)
value NCRYPT_KEY_PROTECTION_INTERFACE (0x00010004)
value NCRYPT_KEY_STORAGE_INTERFACE (0x00010001)
value NCRYPT_MACHINE_KEY_FLAG (0x00000020)
value NCRYPT_MAX_ALG_ID_LENGTH (512)
value NCRYPT_MAX_KEY_NAME_LENGTH (512)
value NCRYPT_MAX_PROPERTY_DATA (0x100000)
value NCRYPT_MAX_PROPERTY_NAME (64)
value NCRYPT_NO_CACHED_PASSWORD (0x00004000)
value NCRYPT_NO_KEY_VALIDATION (BCRYPT_NO_KEY_VALIDATION)
value NCRYPT_NO_PADDING_FLAG (0x00000001)
value NCRYPT_OVERWRITE_KEY_FLAG (0x00000080)
value NCRYPT_PAD_CIPHER_FLAG (0x00000010)
value NCRYPT_PAD_OAEP_FLAG (0x00000004)
value NCRYPT_PAD_PSS_FLAG (0x00000008)
value NCRYPT_PCP_ENCRYPTION_KEY ((0x00000002))
value NCRYPT_PCP_GENERIC_KEY ((NCRYPT_PCP_SIGNATURE_KEY | NCRYPT_PCP_ENCRYPTION_KEY))
value NCRYPT_PCP_HMACVERIFICATION_KEY ((0x00000010))
value NCRYPT_PCP_IDENTITY_KEY ((0x00000008))
value NCRYPT_PCP_SIGNATURE_KEY ((0x00000001))
value NCRYPT_PCP_STORAGE_KEY ((0x00000004))
value NCRYPT_PERSIST_FLAG (0x80000000)
value NCRYPT_PERSIST_ONLY_FLAG (0x40000000)
value NCRYPT_PIN_CACHE_APPLICATION_TICKET_BYTE_LENGTH (90)
value NCRYPT_PIN_CACHE_CLEAR_FOR_CALLING_PROCESS_OPTION (0x00000001)
value NCRYPT_PIN_CACHE_DISABLE_DPL_FLAG (0x00000001)
value NCRYPT_PIN_CACHE_PIN_BYTE_LENGTH (90)
value NCRYPT_PIN_CACHE_REQUIRE_GESTURE_FLAG (0x00000001)
value NCRYPT_PLATFORM_ATTEST_MAGIC (0x44504150)
value NCRYPT_PREFER_VIRTUAL_ISOLATION_FLAG (0x00010000)
value NCRYPT_PROTECTED_KEY_BLOB_MAGIC (0x4B545250)
value NCRYPT_PROTECT_TO_LOCAL_SYSTEM (0x00008000)
value NCRYPT_PUBLIC_LENGTH_PROPERTY (BCRYPT_PUBLIC_KEY_LENGTH)
value NCRYPT_REGISTER_NOTIFY_FLAG (0x00000001)
value NCRYPT_RNG_OPERATION (BCRYPT_RNG_OPERATION)
value NCRYPT_RSA_ALGORITHM (BCRYPT_RSA_ALGORITHM)
value NCRYPT_RSA_ALGORITHM_GROUP (NCRYPT_RSA_ALGORITHM)
value NCRYPT_RSA_SIGN_ALGORITHM (BCRYPT_RSA_SIGN_ALGORITHM)
value NCRYPT_SCHANNEL_INTERFACE (0x00010002)
value NCRYPT_SCHANNEL_SIGNATURE_INTERFACE (0x00010003)
value NCRYPT_SEALING_FLAG (0x00000100)
value NCRYPT_SECRET_AGREEMENT_INTERFACE (BCRYPT_SECRET_AGREEMENT_INTERFACE)
value NCRYPT_SECRET_AGREEMENT_OPERATION (BCRYPT_SECRET_AGREEMENT_OPERATION)
value NCRYPT_SIGNATURE_INTERFACE (BCRYPT_SIGNATURE_INTERFACE)
value NCRYPT_SIGNATURE_LENGTH_PROPERTY (BCRYPT_SIGNATURE_LENGTH)
value NCRYPT_SIGNATURE_OPERATION (BCRYPT_SIGNATURE_OPERATION)
value NCRYPT_SILENT_FLAG (0x00000040)
value NCRYPT_TPM_LOADABLE_KEY_BLOB_MAGIC (0x4D54504B)
value NCRYPT_TPM_PAD_PSS_IGNORE_SALT (0x00000020)
value NCRYPT_TPM_PLATFORM_ATTESTATION_STATEMENT_CURRENT_VERSION (NCRYPT_TPM_PLATFORM_ATTESTATION_STATEMENT_V0)
value NCRYPT_TPM_PSS_SALT_SIZE_HASHSIZE (0x00000002)
value NCRYPT_TPM_PSS_SALT_SIZE_MAXIMUM (0x00000001)
value NCRYPT_TPM_PSS_SALT_SIZE_UNKNOWN (0x00000000)
value NCRYPT_TREAT_NIST_AS_GENERIC_ECC_FLAG (0x00002000)
value NCRYPT_UI_APPCONTAINER_ACCESS_MEDIUM_FLAG (0x00000008)
value NCRYPT_UI_FINGERPRINT_PROTECTION_FLAG (0x00000004)
value NCRYPT_UI_FORCE_HIGH_PROTECTION_FLAG (0x00000002)
value NCRYPT_UI_PROTECT_KEY_FLAG (0x00000001)
value NCRYPT_UNREGISTER_NOTIFY_FLAG (0x00000002)
value NCRYPT_USE_PER_BOOT_KEY_FLAG (0x00040000)
value NCRYPT_USE_VIRTUAL_ISOLATION_FLAG (0x00020000)
value NCRYPT_VSM_KEY_ATTESTATION_CLAIM_RESTRICTIONS_CURRENT_VERSION (NCRYPT_VSM_KEY_ATTESTATION_CLAIM_RESTRICTIONS_V0)
value NCRYPT_VSM_KEY_ATTESTATION_STATEMENT_CURRENT_VERSION (NCRYPT_VSM_KEY_ATTESTATION_STATEMENT_V0)
value NCRYPT_WRITE_KEY_TO_LEGACY_STORE_FLAG (0x00000200)
value NDR_CUSTOM_OR_DEFAULT_ALLOCATOR (0x10000000UL)
value NDR_DEFAULT_ALLOCATOR (0x20000000UL)
value NDR_LOCAL_ENDIAN (NDR_LITTLE_ENDIAN)
value NETINFO_DISKRED (0x00000004)
value NETINFO_PRINTERRED (0x00000008)
value NETPROPERTY_PERSISTENT (1)
value NETSCAPE_SIGN_CA_CERT_TYPE (0x01)
value NETSCAPE_SIGN_CERT_TYPE (0x10)
value NETSCAPE_SMIME_CA_CERT_TYPE (0x02)
value NETSCAPE_SMIME_CERT_TYPE (0x20)
value NETSCAPE_SSL_CA_CERT_TYPE (0x04)
value NETSCAPE_SSL_CLIENT_AUTH_CERT_TYPE (0x80)
value NETSCAPE_SSL_SERVER_AUTH_CERT_TYPE (0x40)
value NETWORK_APP_INSTANCE_CSV_FLAGS_VALID_ONLY_IF_CSV_COORDINATOR (0x00000001)
value NEWFILEOPENORD (1547)
value NEWFORMATDLGWITHLINK (1591)
value NEWFRAME (1)
value NEWTRANSPARENT (3)
value NEXTBAND (3)
value NFR_ANSI (1)
value NFR_UNICODE (2)
value NF_QUERY (3)
value NF_REQUERY (4)
value NID_EXTERNAL_PEN (0x00000008)
value NID_EXTERNAL_TOUCH (0x00000002)
value NID_INTEGRATED_PEN (0x00000004)
value NID_INTEGRATED_TOUCH (0x00000001)
value NID_MULTI_INPUT (0x00000040)
value NID_READY (0x00000080)
value NIF_GUID (0x00000020)
value NIF_ICON (0x00000002)
value NIF_INFO (0x00000010)
value NIF_MESSAGE (0x00000001)
value NIF_REALTIME (0x00000040)
value NIF_SHOWTIP (0x00000080)
value NIF_STATE (0x00000008)
value NIF_TIP (0x00000004)
value NIIF_ERROR (0x00000003)
value NIIF_ICON_MASK (0x0000000F)
value NIIF_INFO (0x00000001)
value NIIF_LARGE_ICON (0x00000020)
value NIIF_NONE (0x00000000)
value NIIF_NOSOUND (0x00000010)
value NIIF_RESPECT_QUIET_TIME (0x00000080)
value NIIF_USER (0x00000004)
value NIIF_WARNING (0x00000002)
value NIM_ADD (0x00000000)
value NIM_DELETE (0x00000002)
value NIM_MODIFY (0x00000001)
value NIM_SETFOCUS (0x00000003)
value NIM_SETVERSION (0x00000004)
value NINF_KEY (0x1)
value NIN_BALLOONHIDE ((WM_USER + 3))
value NIN_BALLOONSHOW ((WM_USER + 2))
value NIN_BALLOONTIMEOUT ((WM_USER + 4))
value NIN_BALLOONUSERCLICK ((WM_USER + 5))
value NIN_KEYSELECT ((NIN_SELECT | NINF_KEY))
value NIN_POPUPCLOSE ((WM_USER + 7))
value NIN_POPUPOPEN ((WM_USER + 6))
value NIN_SELECT ((WM_USER + 0))
value NIS_HIDDEN (0x00000001)
value NIS_SHAREDICON (0x00000002)
value NI_CHANGECANDIDATELIST (0x0013)
value NI_CLOSECANDIDATE (0x0011)
value NI_COMPOSITIONSTR (0x0015)
value NI_DGRAM (0x10)
value NI_FINALIZECONVERSIONRESULT (0x0014)
value NI_IMEMENUSELECTED (0x0018)
value NI_MAXHOST (1025)
value NI_MAXSERV (32)
value NI_NAMEREQD (0x04)
value NI_NOFQDN (0x01)
value NI_NUMERICHOST (0x02)
value NI_NUMERICSERV (0x08)
value NI_OPENCANDIDATE (0x0010)
value NI_SELECTCANDIDATESTR (0x0012)
value NI_SETCANDIDATE_PAGESIZE (0x0017)
value NI_SETCANDIDATE_PAGESTART (0x0016)
value NLS_ALPHANUMERIC (0x00000000)
value NLS_DBCSCHAR (0x00010000)
value NLS_HIRAGANA (0x00040000)
value NLS_IME_CONVERSION (0x00800000)
value NLS_IME_DISABLE (0x20000000)
value NLS_KATAKANA (0x00020000)
value NLS_ROMAN (0x00400000)
value NLS_VALID_LOCALE_MASK (0x000fffff)
value NMPWAIT_NOWAIT (0x00000001)
value NMPWAIT_USE_DEFAULT_WAIT (0x00000000)
value NMPWAIT_WAIT_FOREVER (0xffffffff)
value NOERROR (0)
value NOMIRRORBITMAP ((DWORD)0x80000000)
value NONANTIALIASED_QUALITY (3)
value NONZEROLHND ((LMEM_MOVEABLE))
value NONZEROLPTR ((LMEM_FIXED))
value NON_PAGED_DEBUG_SIGNATURE (0x494E)
value NOPARITY (0)
value NORMAL_PRINT (( 0x00000000 ))
value NORMAL_PRIORITY_CLASS (0x00000020)
value NORM_IGNORECASE (0x00000001)
value NORM_IGNOREKANATYPE (0x00010000)
value NORM_IGNORENONSPACE (0x00000002)
value NORM_IGNORESYMBOLS (0x00000004)
value NORM_IGNOREWIDTH (0x00020000)
value NORM_LINGUISTIC_CASING (0x08000000)
value NOTIFYICON_VERSION (3)
value NOTSRCCOPY ((DWORD)0x00330008)
value NOTSRCERASE ((DWORD)0x001100A6)
value NO_ADDRESS (WSANO_ADDRESS)
value NO_DATA (WSANO_DATA)
value NO_ERROR (0)
value NO_PRIORITY (0)
value NO_PROPAGATE_INHERIT_ACE ((0x4))
value NO_RECOVERY (WSANO_RECOVERY)
value NRC_ACTSES (0x0f)
value NRC_BADDR (0x07)
value NRC_BRIDGE (0x23)
value NRC_BUFLEN (0x01)
value NRC_CANCEL (0x26)
value NRC_CANOCCR (0x24)
value NRC_CMDCAN (0x0b)
value NRC_CMDTMO (0x05)
value NRC_DUPENV (0x30)
value NRC_DUPNAME (0x0d)
value NRC_ENVNOTDEF (0x34)
value NRC_GOODRET (0x00)
value NRC_IFBUSY (0x21)
value NRC_ILLCMD (0x03)
value NRC_ILLNN (0x13)
value NRC_INCOMP (0x06)
value NRC_INUSE (0x16)
value NRC_INVADDRESS (0x39)
value NRC_INVDDID (0x3B)
value NRC_LOCKFAIL (0x3C)
value NRC_LOCTFUL (0x11)
value NRC_MAXAPPS (0x36)
value NRC_NAMCONF (0x19)
value NRC_NAMERR (0x17)
value NRC_NAMTFUL (0x0e)
value NRC_NOCALL (0x14)
value NRC_NORES (0x09)
value NRC_NORESOURCES (0x38)
value NRC_NOSAPS (0x37)
value NRC_NOWILD (0x15)
value NRC_OPENERR (0x3f)
value NRC_OSRESNOTAV (0x35)
value NRC_PENDING (0xff)
value NRC_REMTFUL (0x12)
value NRC_SABORT (0x18)
value NRC_SCLOSED (0x0a)
value NRC_SNUMOUT (0x08)
value NRC_SYSTEM (0x40)
value NRC_TOOMANY (0x22)
value NS_ALL ((0))
value NS_BTH ((16))
value NS_DHCP ((6))
value NS_DNS ((12))
value NS_EMAIL ((37))
value NS_LOCALNAME ((19))
value NS_MS ((30))
value NS_NBP ((20))
value NS_NDS ((2))
value NS_NETBT ((13))
value NS_NETDES ((60))
value NS_NIS ((41))
value NS_NISPLUS ((42))
value NS_NLA ((15))
value NS_NTDS ((32))
value NS_PEER_BROWSE ((3))
value NS_PNRPCLOUD ((39))
value NS_PNRPNAME ((38))
value NS_SAP ((1))
value NS_SLP ((5))
value NS_STDA ((31))
value NS_TCPIP_HOSTS ((11))
value NS_TCPIP_LOCAL ((10))
value NS_WINS ((14))
value NS_WRQ ((50))
value NTAPI_INLINE (NTAPI)
value NTDDI_LONGHORN (NTDDI_VISTA)
value NTDDI_VERSION (WDK_NTDDI_VERSION)
value NTDDI_VISTA (NTDDI_WIN6)
value NTDDI_WINBLUE (0x06030000)
value NTDDI_WINTHRESHOLD (0x0A000000)
value NTDDI_WINXP (0x05010000)
value NTE_AUTHENTICATION_IGNORED (_HRESULT_TYPEDEF_(0x80090031L))
value NTE_BAD_ALGID (_HRESULT_TYPEDEF_(0x80090008L))
value NTE_BAD_DATA (_HRESULT_TYPEDEF_(0x80090005L))
value NTE_BAD_FLAGS (_HRESULT_TYPEDEF_(0x80090009L))
value NTE_BAD_HASH (_HRESULT_TYPEDEF_(0x80090002L))
value NTE_BAD_HASH_STATE (_HRESULT_TYPEDEF_(0x8009000CL))
value NTE_BAD_KEY (_HRESULT_TYPEDEF_(0x80090003L))
value NTE_BAD_KEYSET (_HRESULT_TYPEDEF_(0x80090016L))
value NTE_BAD_KEYSET_PARAM (_HRESULT_TYPEDEF_(0x8009001FL))
value NTE_BAD_KEY_STATE (_HRESULT_TYPEDEF_(0x8009000BL))
value NTE_BAD_LEN (_HRESULT_TYPEDEF_(0x80090004L))
value NTE_BAD_PROVIDER (_HRESULT_TYPEDEF_(0x80090013L))
value NTE_BAD_PROV_TYPE (_HRESULT_TYPEDEF_(0x80090014L))
value NTE_BAD_PUBLIC_KEY (_HRESULT_TYPEDEF_(0x80090015L))
value NTE_BAD_SIGNATURE (_HRESULT_TYPEDEF_(0x80090006L))
value NTE_BAD_TYPE (_HRESULT_TYPEDEF_(0x8009000AL))
value NTE_BAD_UID (_HRESULT_TYPEDEF_(0x80090001L))
value NTE_BAD_VER (_HRESULT_TYPEDEF_(0x80090007L))
value NTE_BUFFERS_OVERLAP (_HRESULT_TYPEDEF_(0x8009002BL))
value NTE_BUFFER_TOO_SMALL (_HRESULT_TYPEDEF_(0x80090028L))
value NTE_DECRYPTION_FAILURE (_HRESULT_TYPEDEF_(0x8009002CL))
value NTE_DEVICE_NOT_FOUND (_HRESULT_TYPEDEF_(0x80090035L))
value NTE_DEVICE_NOT_READY (_HRESULT_TYPEDEF_(0x80090030L))
value NTE_DOUBLE_ENCRYPT (_HRESULT_TYPEDEF_(0x80090012L))
value NTE_ENCRYPTION_FAILURE (_HRESULT_TYPEDEF_(0x80090034L))
value NTE_EXISTS (_HRESULT_TYPEDEF_(0x8009000FL))
value NTE_FAIL (_HRESULT_TYPEDEF_(0x80090020L))
value NTE_FIXEDPARAMETER (_HRESULT_TYPEDEF_(0x80090025L))
value NTE_HMAC_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8009002FL))
value NTE_INCORRECT_PASSWORD (_HRESULT_TYPEDEF_(0x80090033L))
value NTE_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x8009002DL))
value NTE_INVALID_HANDLE (_HRESULT_TYPEDEF_(0x80090026L))
value NTE_INVALID_PARAMETER (_HRESULT_TYPEDEF_(0x80090027L))
value NTE_KEYSET_ENTRY_BAD (_HRESULT_TYPEDEF_(0x8009001AL))
value NTE_KEYSET_NOT_DEF (_HRESULT_TYPEDEF_(0x80090019L))
value NTE_NOT_ACTIVE_CONSOLE (_HRESULT_TYPEDEF_(0x80090038L))
value NTE_NOT_FOUND (_HRESULT_TYPEDEF_(0x80090011L))
value NTE_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80090029L))
value NTE_NO_KEY (_HRESULT_TYPEDEF_(0x8009000DL))
value NTE_NO_MEMORY (_HRESULT_TYPEDEF_(0x8009000EL))
value NTE_NO_MORE_ITEMS (_HRESULT_TYPEDEF_(0x8009002AL))
value NTE_OP_OK (0)
value NTE_PASSWORD_CHANGE_REQUIRED (_HRESULT_TYPEDEF_(0x80090037L))
value NTE_PERM (_HRESULT_TYPEDEF_(0x80090010L))
value NTE_PROVIDER_DLL_FAIL (_HRESULT_TYPEDEF_(0x8009001DL))
value NTE_PROV_DLL_NOT_FOUND (_HRESULT_TYPEDEF_(0x8009001EL))
value NTE_PROV_TYPE_ENTRY_BAD (_HRESULT_TYPEDEF_(0x80090018L))
value NTE_PROV_TYPE_NOT_DEF (_HRESULT_TYPEDEF_(0x80090017L))
value NTE_PROV_TYPE_NO_MATCH (_HRESULT_TYPEDEF_(0x8009001BL))
value NTE_SIGNATURE_FILE_BAD (_HRESULT_TYPEDEF_(0x8009001CL))
value NTE_SILENT_CONTEXT (_HRESULT_TYPEDEF_(0x80090022L))
value NTE_SYS_ERR (_HRESULT_TYPEDEF_(0x80090021L))
value NTE_TEMPORARY_PROFILE (_HRESULT_TYPEDEF_(0x80090024L))
value NTE_TOKEN_KEYSET_STORAGE_FULL (_HRESULT_TYPEDEF_(0x80090023L))
value NTE_UI_REQUIRED (_HRESULT_TYPEDEF_(0x8009002EL))
value NTE_USER_CANCELLED (_HRESULT_TYPEDEF_(0x80090036L))
value NTE_VALIDATION_FAILED (_HRESULT_TYPEDEF_(0x80090032L))
value NTM_BOLD (0x00000020L)
value NTM_DSIG (0x00200000)
value NTM_ITALIC (0x00000001L)
value NTM_MULTIPLEMASTER (0x00080000)
value NTM_NONNEGATIVE_AC (0x00010000)
value NTM_PS_OPENTYPE (0x00020000)
value NTM_REGULAR (0x00000040L)
value NTM_TT_OPENTYPE (0x00040000)
value NTSYSAPI (DECLSPEC_IMPORT)
value NTSYSCALLAPI (DECLSPEC_IMPORT)
value NULLREGION (1)
value NULL_BRUSH (5)
value NULL_PEN (8)
value NUMA_NO_PREFERRED_NODE (((DWORD) -1))
value NUMBRUSHES (16)
value NUMCOLORS (24)
value NUMFONTS (22)
value NUMLOCK_ON (0x0020)
value NUMMARKERS (20)
value NUMPENS (18)
value NUMPRS_CURRENCY (0x0400)
value NUMPRS_DECIMAL (0x0100)
value NUMPRS_EXPONENT (0x0800)
value NUMPRS_HEX_OCT (0x0040)
value NUMPRS_INEXACT (0x20000)
value NUMPRS_LEADING_MINUS (0x0010)
value NUMPRS_LEADING_PLUS (0x0004)
value NUMPRS_LEADING_WHITE (0x0001)
value NUMPRS_NEG (0x10000)
value NUMPRS_PARENS (0x0080)
value NUMPRS_STD (0x1FFF)
value NUMPRS_THOUSANDS (0x0200)
value NUMPRS_TRAILING_MINUS (0x0020)
value NUMPRS_TRAILING_PLUS (0x0008)
value NUMPRS_TRAILING_WHITE (0x0002)
value NUMPRS_USE_ALL (0x1000)
value NUMRESERVED (106)
value NUM_DISCHARGE_POLICIES (4)
value N_BTMASK (0x000F)
value N_BTSHFT (4)
value N_TMASK (0x0030)
value N_TSHIFT (2)
value OBJECT_INHERIT_ACE ((0x1))
value OBJID_ALERT (((LONG)0xFFFFFFF6))
value OBJID_CARET (((LONG)0xFFFFFFF8))
value OBJID_CLIENT (((LONG)0xFFFFFFFC))
value OBJID_CURSOR (((LONG)0xFFFFFFF7))
value OBJID_HSCROLL (((LONG)0xFFFFFFFA))
value OBJID_MENU (((LONG)0xFFFFFFFD))
value OBJID_NATIVEOM (((LONG)0xFFFFFFF0))
value OBJID_QUERYCLASSNAMEIDX (((LONG)0xFFFFFFF4))
value OBJID_SIZEGRIP (((LONG)0xFFFFFFF9))
value OBJID_SOUND (((LONG)0xFFFFFFF5))
value OBJID_SYSMENU (((LONG)0xFFFFFFFF))
value OBJID_TITLEBAR (((LONG)0xFFFFFFFE))
value OBJID_VSCROLL (((LONG)0xFFFFFFFB))
value OBJID_WINDOW (((LONG)0x00000000))
value OBJ_BITMAP (7)
value OBJ_BRUSH (2)
value OBJ_COLORSPACE (14)
value OBJ_DC (3)
value OBJ_ENHMETADC (12)
value OBJ_ENHMETAFILE (13)
value OBJ_EXTPEN (11)
value OBJ_FONT (6)
value OBJ_MEMDC (10)
value OBJ_METADC (4)
value OBJ_METAFILE (9)
value OBJ_PAL (5)
value OBJ_PEN (1)
value OBJ_REGION (8)
value OCSP_BASIC_BY_KEY_RESPONDER_ID (2)
value OCSP_BASIC_BY_NAME_RESPONDER_ID (1)
value OCSP_BASIC_GOOD_CERT_STATUS (0)
value OCSP_BASIC_RESPONSE (((LPCSTR) 69))
value OCSP_BASIC_REVOKED_CERT_STATUS (1)
value OCSP_BASIC_SIGNED_RESPONSE (((LPCSTR) 68))
value OCSP_BASIC_UNKNOWN_CERT_STATUS (2)
value OCSP_INTERNAL_ERROR_RESPONSE (2)
value OCSP_MALFORMED_REQUEST_RESPONSE (1)
value OCSP_REQUEST (((LPCSTR) 66))
value OCSP_RESPONSE (((LPCSTR) 67))
value OCSP_SIGNED_REQUEST (((LPCSTR) 65))
value OCSP_SIG_REQUIRED_RESPONSE (5)
value OCSP_SUCCESSFUL_RESPONSE (0)
value OCSP_TRY_LATER_RESPONSE (3)
value OCSP_UNAUTHORIZED_RESPONSE (6)
value ODA_DRAWENTIRE (0x0001)
value ODA_FOCUS (0x0004)
value ODA_SELECT (0x0002)
value ODDPARITY (1)
value ODS_CHECKED (0x0008)
value ODS_COMBOBOXEDIT (0x1000)
value ODS_DEFAULT (0x0020)
value ODS_DISABLED (0x0004)
value ODS_FOCUS (0x0010)
value ODS_GRAYED (0x0002)
value ODS_HOTLIGHT (0x0040)
value ODS_INACTIVE (0x0080)
value ODS_NOACCEL (0x0100)
value ODS_NOFOCUSRECT (0x0200)
value ODS_SELECTED (0x0001)
value ODT_BUTTON (4)
value ODT_COMBOBOX (3)
value ODT_LISTBOX (2)
value ODT_MENU (1)
value ODT_STATIC (5)
value OEM_CHARSET (255)
value OEM_FIXED_FONT (10)
value OFFLINE_STATUS_INCOMPLETE (0x0004)
value OFFLINE_STATUS_LOCAL (0x0001)
value OFFLINE_STATUS_REMOTE (0x0002)
value OFFLOAD_READ_FLAG_ALL_ZERO_BEYOND_CURRENT_RANGE ((1))
value OFN_ALLOWMULTISELECT (0x00000200)
value OFN_CREATEPROMPT (0x00002000)
value OFN_DONTADDTORECENT (0x02000000)
value OFN_ENABLEHOOK (0x00000020)
value OFN_ENABLEINCLUDENOTIFY (0x00400000)
value OFN_ENABLESIZING (0x00800000)
value OFN_ENABLETEMPLATE (0x00000040)
value OFN_ENABLETEMPLATEHANDLE (0x00000080)
value OFN_EXPLORER (0x00080000)
value OFN_EXTENSIONDIFFERENT (0x00000400)
value OFN_EX_NOPLACESBAR (0x00000001)
value OFN_FILEMUSTEXIST (0x00001000)
value OFN_FORCESHOWHIDDEN (0x10000000)
value OFN_HIDEREADONLY (0x00000004)
value OFN_LONGNAMES (0x00200000)
value OFN_NOCHANGEDIR (0x00000008)
value OFN_NODEREFERENCELINKS (0x00100000)
value OFN_NOLONGNAMES (0x00040000)
value OFN_NONETWORKBUTTON (0x00020000)
value OFN_NOREADONLYRETURN (0x00008000)
value OFN_NOTESTFILECREATE (0x00010000)
value OFN_NOVALIDATE (0x00000100)
value OFN_OVERWRITEPROMPT (0x00000002)
value OFN_PATHMUSTEXIST (0x00000800)
value OFN_READONLY (0x00000001)
value OFN_SHAREAWARE (0x00004000)
value OFN_SHAREFALLTHROUGH (2)
value OFN_SHARENOWARN (1)
value OFN_SHAREWARN (0)
value OFN_SHOWHELP (0x00000010)
value OFS_MAXPATHNAME (128)
value OF_CANCEL (0x00000800)
value OF_CREATE (0x00001000)
value OF_DELETE (0x00000200)
value OF_EXIST (0x00004000)
value OF_PARSE (0x00000100)
value OF_PROMPT (0x00002000)
value OF_READ (0x00000000)
value OF_READWRITE (0x00000002)
value OF_REOPEN (0x00008000)
value OF_SHARE_COMPAT (0x00000000)
value OF_SHARE_DENY_NONE (0x00000040)
value OF_SHARE_DENY_READ (0x00000030)
value OF_SHARE_DENY_WRITE (0x00000020)
value OF_SHARE_EXCLUSIVE (0x00000010)
value OF_VERIFY (0x00000400)
value OF_WRITE (0x00000001)
value OLDFONTENUMPROC (OLDFONTENUMPROCA)
value OLECREATE_LEAVERUNNING (0x00000001)
value OLEIVERB_DISCARDUNDOSTATE ((-6L))
value OLEIVERB_HIDE ((-3L))
value OLEIVERB_INPLACEACTIVATE ((-5L))
value OLEIVERB_OPEN ((-2L))
value OLEIVERB_PRIMARY ((0L))
value OLEIVERB_SHOW ((-1L))
value OLEIVERB_UIACTIVATE ((-4L))
value OLEOBJ_E_FIRST (0x80040180L)
value OLEOBJ_E_INVALIDVERB (_HRESULT_TYPEDEF_(0x80040181L))
value OLEOBJ_E_LAST (0x8004018FL)
value OLEOBJ_E_NOVERBS (_HRESULT_TYPEDEF_(0x80040180L))
value OLEOBJ_S_CANNOT_DOVERB_NOW (_HRESULT_TYPEDEF_(0x00040181L))
value OLEOBJ_S_FIRST (0x00040180L)
value OLEOBJ_S_INVALIDHWND (_HRESULT_TYPEDEF_(0x00040182L))
value OLEOBJ_S_INVALIDVERB (_HRESULT_TYPEDEF_(0x00040180L))
value OLEOBJ_S_LAST (0x0004018FL)
value OLE_E_ADVF (_HRESULT_TYPEDEF_(0x80040001L))
value OLE_E_ADVISENOTSUPPORTED (_HRESULT_TYPEDEF_(0x80040003L))
value OLE_E_BLANK (_HRESULT_TYPEDEF_(0x80040007L))
value OLE_E_CANTCONVERT (_HRESULT_TYPEDEF_(0x80040011L))
value OLE_E_CANT_BINDTOSOURCE (_HRESULT_TYPEDEF_(0x8004000AL))
value OLE_E_CANT_GETMONIKER (_HRESULT_TYPEDEF_(0x80040009L))
value OLE_E_CLASSDIFF (_HRESULT_TYPEDEF_(0x80040008L))
value OLE_E_ENUM_NOMORE (_HRESULT_TYPEDEF_(0x80040002L))
value OLE_E_FIRST (((HRESULT)0x80040000L))
value OLE_E_INVALIDHWND (_HRESULT_TYPEDEF_(0x8004000FL))
value OLE_E_INVALIDRECT (_HRESULT_TYPEDEF_(0x8004000DL))
value OLE_E_LAST (((HRESULT)0x800400FFL))
value OLE_E_NOCACHE (_HRESULT_TYPEDEF_(0x80040006L))
value OLE_E_NOCONNECTION (_HRESULT_TYPEDEF_(0x80040004L))
value OLE_E_NOSTORAGE (_HRESULT_TYPEDEF_(0x80040012L))
value OLE_E_NOTRUNNING (_HRESULT_TYPEDEF_(0x80040005L))
value OLE_E_NOT_INPLACEACTIVE (_HRESULT_TYPEDEF_(0x80040010L))
value OLE_E_OLEVERB (_HRESULT_TYPEDEF_(0x80040000L))
value OLE_E_PROMPTSAVECANCELLED (_HRESULT_TYPEDEF_(0x8004000CL))
value OLE_E_STATIC (_HRESULT_TYPEDEF_(0x8004000BL))
value OLE_E_WRONGCOMPOBJ (_HRESULT_TYPEDEF_(0x8004000EL))
value OLE_S_FIRST (((HRESULT)0x00040000L))
value OLE_S_LAST (((HRESULT)0x000400FFL))
value OLE_S_MAC_CLIPFORMAT (_HRESULT_TYPEDEF_(0x00040002L))
value OLE_S_STATIC (_HRESULT_TYPEDEF_(0x00040001L))
value OLE_S_USEREG (_HRESULT_TYPEDEF_(0x00040000L))
value ONESTOPBIT (0)
value ONL_CONNECTION_COUNT_LIMIT (_HRESULT_TYPEDEF_(0x8086000DL))
value ONL_E_ACCESS_DENIED_BY_TOU (_HRESULT_TYPEDEF_(0x80860002L))
value ONL_E_ACCOUNT_LOCKED (_HRESULT_TYPEDEF_(0x80860007L))
value ONL_E_ACCOUNT_SUSPENDED_ABUSE (_HRESULT_TYPEDEF_(0x8086000BL))
value ONL_E_ACCOUNT_SUSPENDED_COMPROIMISE (_HRESULT_TYPEDEF_(0x8086000AL))
value ONL_E_ACCOUNT_UPDATE_REQUIRED (_HRESULT_TYPEDEF_(0x80860005L))
value ONL_E_ACTION_REQUIRED (_HRESULT_TYPEDEF_(0x8086000CL))
value ONL_E_CONNECTED_ACCOUNT_CAN_NOT_SIGNOUT (_HRESULT_TYPEDEF_(0x8086000EL))
value ONL_E_EMAIL_VERIFICATION_REQUIRED (_HRESULT_TYPEDEF_(0x80860009L))
value ONL_E_FORCESIGNIN (_HRESULT_TYPEDEF_(0x80860006L))
value ONL_E_INVALID_APPLICATION (_HRESULT_TYPEDEF_(0x80860003L))
value ONL_E_INVALID_AUTHENTICATION_TARGET (_HRESULT_TYPEDEF_(0x80860001L))
value ONL_E_PARENTAL_CONSENT_REQUIRED (_HRESULT_TYPEDEF_(0x80860008L))
value ONL_E_PASSWORD_UPDATE_REQUIRED (_HRESULT_TYPEDEF_(0x80860004L))
value ONL_E_REQUEST_THROTTLED (_HRESULT_TYPEDEF_(0x80860010L))
value ONL_E_USER_AUTHENTICATION_REQUIRED (_HRESULT_TYPEDEF_(0x8086000FL))
value OPAQUE (2)
value OPAQUEKEYBLOB (0x9)
value OPENCARDNAMEA_EX (OPENCARDNAME_EXA)
value OPENCARDNAMEW_EX (OPENCARDNAME_EXW)
value OPENCARDNAME_A (OPENCARDNAMEA)
value OPENCARDNAME_W (OPENCARDNAMEW)
value OPENCHANNEL (4110)
value OPEN_ALWAYS (4)
value OPEN_EXISTING (3)
value OPERATION_API_VERSION (1)
value OPERATION_END_DISCARD (0x1)
value OPERATION_START_TRACE_CURRENT_THREAD (0x1)
value OPLOCK_LEVEL_CACHE_HANDLE ((0x00000002))
value OPLOCK_LEVEL_CACHE_READ ((0x00000001))
value OPLOCK_LEVEL_CACHE_WRITE ((0x00000004))
value ORD_LANGDRIVER (1)
value OR_INVALID_OID (1911)
value OR_INVALID_OXID (1910)
value OR_INVALID_SET (1912)
value OSS_ACCESS_SERIALIZATION_ERROR (_HRESULT_TYPEDEF_(0x80093013L))
value OSS_API_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x80093029L))
value OSS_BAD_ARG (_HRESULT_TYPEDEF_(0x80093006L))
value OSS_BAD_ENCRULES (_HRESULT_TYPEDEF_(0x80093016L))
value OSS_BAD_PTR (_HRESULT_TYPEDEF_(0x8009300BL))
value OSS_BAD_TABLE (_HRESULT_TYPEDEF_(0x8009300FL))
value OSS_BAD_TIME (_HRESULT_TYPEDEF_(0x8009300CL))
value OSS_BAD_VERSION (_HRESULT_TYPEDEF_(0x80093007L))
value OSS_BERDER_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x8009302AL))
value OSS_CANT_CLOSE_TRACE_FILE (_HRESULT_TYPEDEF_(0x8009302EL))
value OSS_CANT_OPEN_TRACE_FILE (_HRESULT_TYPEDEF_(0x8009301BL))
value OSS_CANT_OPEN_TRACE_WINDOW (_HRESULT_TYPEDEF_(0x80093018L))
value OSS_COMPARATOR_CODE_NOT_LINKED (_HRESULT_TYPEDEF_(0x80093025L))
value OSS_COMPARATOR_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x80093024L))
value OSS_CONSTRAINT_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x80093023L))
value OSS_CONSTRAINT_VIOLATED (_HRESULT_TYPEDEF_(0x80093011L))
value OSS_COPIER_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x80093022L))
value OSS_DATA_ERROR (_HRESULT_TYPEDEF_(0x80093005L))
value OSS_FATAL_ERROR (_HRESULT_TYPEDEF_(0x80093012L))
value OSS_INDEFINITE_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8009300DL))
value OSS_LIMITED (_HRESULT_TYPEDEF_(0x8009300AL))
value OSS_MEM_ERROR (_HRESULT_TYPEDEF_(0x8009300EL))
value OSS_MEM_MGR_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x80093026L))
value OSS_MORE_BUF (_HRESULT_TYPEDEF_(0x80093001L))
value OSS_MORE_INPUT (_HRESULT_TYPEDEF_(0x80093004L))
value OSS_MUTEX_NOT_CREATED (_HRESULT_TYPEDEF_(0x8009302DL))
value OSS_NEGATIVE_UINTEGER (_HRESULT_TYPEDEF_(0x80093002L))
value OSS_NULL_FCN (_HRESULT_TYPEDEF_(0x80093015L))
value OSS_NULL_TBL (_HRESULT_TYPEDEF_(0x80093014L))
value OSS_OID_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x8009301AL))
value OSS_OPEN_TYPE_ERROR (_HRESULT_TYPEDEF_(0x8009302CL))
value OSS_OUT_MEMORY (_HRESULT_TYPEDEF_(0x80093008L))
value OSS_OUT_OF_RANGE (_HRESULT_TYPEDEF_(0x80093021L))
value OSS_PDU_MISMATCH (_HRESULT_TYPEDEF_(0x80093009L))
value OSS_PDU_RANGE (_HRESULT_TYPEDEF_(0x80093003L))
value OSS_PDV_CODE_NOT_LINKED (_HRESULT_TYPEDEF_(0x80093028L))
value OSS_PDV_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x80093027L))
value OSS_PER_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x8009302BL))
value OSS_REAL_CODE_NOT_LINKED (_HRESULT_TYPEDEF_(0x80093020L))
value OSS_REAL_DLL_NOT_LINKED (_HRESULT_TYPEDEF_(0x8009301FL))
value OSS_TABLE_MISMATCH (_HRESULT_TYPEDEF_(0x8009301DL))
value OSS_TOO_LONG (_HRESULT_TYPEDEF_(0x80093010L))
value OSS_TRACE_FILE_ALREADY_OPEN (_HRESULT_TYPEDEF_(0x8009301CL))
value OSS_TYPE_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8009301EL))
value OSS_UNAVAIL_ENCRULES (_HRESULT_TYPEDEF_(0x80093017L))
value OSS_UNIMPLEMENTED (_HRESULT_TYPEDEF_(0x80093019L))
value OSVERSION_MASK (0xFFFF0000)
value OUTPUT_DEBUG_STRING_EVENT (8)
value OUT_CHARACTER_PRECIS (2)
value OUT_DEFAULT_PRECIS (0)
value OUT_DEVICE_PRECIS (5)
value OUT_OUTLINE_PRECIS (8)
value OUT_PS_ONLY_PRECIS (10)
value OUT_RASTER_PRECIS (6)
value OUT_SCREEN_OUTLINE_PRECIS (9)
value OUT_STRING_PRECIS (1)
value OUT_STROKE_PRECIS (3)
value OUT_TT_ONLY_PRECIS (7)
value OUT_TT_PRECIS (4)
value OVERWRITE_HIDDEN ((4))
value OWNER_SECURITY_INFORMATION ((0x00000001L))
value O_APPEND (_O_APPEND)
value O_BINARY (_O_BINARY)
value O_CREAT (_O_CREAT)
value O_EXCL (_O_EXCL)
value O_NOINHERIT (_O_NOINHERIT)
value O_RANDOM (_O_RANDOM)
value O_RAW (_O_BINARY)
value O_RDONLY (_O_RDONLY)
value O_RDWR (_O_RDWR)
value O_SEQUENTIAL (_O_SEQUENTIAL)
value O_TEMPORARY (_O_TEMPORARY)
value O_TEXT (_O_TEXT)
value O_TRUNC (_O_TRUNC)
value O_WRONLY (_O_WRONLY)
value PAGESETUPDLGORD (1546)
value PAGESETUPDLGORDMOTIF (1550)
value PAGE_ENCLAVE_DECOMMIT ((PAGE_ENCLAVE_MASK | 0))
value PAGE_ENCLAVE_MASK (0x10000000)
value PAGE_ENCLAVE_SS_FIRST ((PAGE_ENCLAVE_MASK | 1))
value PAGE_ENCLAVE_SS_REST ((PAGE_ENCLAVE_MASK | 2))
value PAGE_ENCLAVE_THREAD_CONTROL (0x80000000)
value PAGE_ENCLAVE_UNVALIDATED (0x20000000)
value PAGE_EXECUTE (0x10)
value PAGE_EXECUTE_READ (0x20)
value PAGE_EXECUTE_READWRITE (0x40)
value PAGE_EXECUTE_WRITECOPY (0x80)
value PAGE_GRAPHICS_COHERENT (0x20000)
value PAGE_GRAPHICS_EXECUTE (0x4000)
value PAGE_GRAPHICS_EXECUTE_READ (0x8000)
value PAGE_GRAPHICS_EXECUTE_READWRITE (0x10000)
value PAGE_GRAPHICS_NOACCESS (0x0800)
value PAGE_GRAPHICS_NOCACHE (0x40000)
value PAGE_GRAPHICS_READONLY (0x1000)
value PAGE_GRAPHICS_READWRITE (0x2000)
value PAGE_GUARD (0x100)
value PAGE_NOACCESS (0x01)
value PAGE_NOCACHE (0x200)
value PAGE_READONLY (0x02)
value PAGE_READWRITE (0x04)
value PAGE_REVERT_TO_FILE_MAP (0x80000000)
value PAGE_TARGETS_INVALID (0x40000000)
value PAGE_TARGETS_NO_UPDATE (0x40000000)
value PAGE_WRITECOMBINE (0x400)
value PAGE_WRITECOPY (0x08)
value PANOSE_COUNT (10)
value PAN_ANY (0)
value PAN_ARMSTYLE_INDEX (6)
value PAN_BENT_ARMS_DOUBLE_SERIF (11)
value PAN_BENT_ARMS_HORZ (7)
value PAN_BENT_ARMS_SINGLE_SERIF (10)
value PAN_BENT_ARMS_VERT (9)
value PAN_BENT_ARMS_WEDGE (8)
value PAN_CONTRAST_HIGH (8)
value PAN_CONTRAST_INDEX (4)
value PAN_CONTRAST_LOW (4)
value PAN_CONTRAST_MEDIUM (6)
value PAN_CONTRAST_MEDIUM_HIGH (7)
value PAN_CONTRAST_MEDIUM_LOW (5)
value PAN_CONTRAST_NONE (2)
value PAN_CONTRAST_VERY_HIGH (9)
value PAN_CONTRAST_VERY_LOW (3)
value PAN_CULTURE_LATIN (0)
value PAN_FAMILYTYPE_INDEX (0)
value PAN_FAMILY_DECORATIVE (4)
value PAN_FAMILY_PICTORIAL (5)
value PAN_FAMILY_SCRIPT (3)
value PAN_FAMILY_TEXT_DISPLAY (2)
value PAN_LETTERFORM_INDEX (7)
value PAN_LETT_NORMAL_BOXED (4)
value PAN_LETT_NORMAL_CONTACT (2)
value PAN_LETT_NORMAL_FLATTENED (5)
value PAN_LETT_NORMAL_OFF_CENTER (7)
value PAN_LETT_NORMAL_ROUNDED (6)
value PAN_LETT_NORMAL_SQUARE (8)
value PAN_LETT_NORMAL_WEIGHTED (3)
value PAN_LETT_OBLIQUE_BOXED (11)
value PAN_LETT_OBLIQUE_CONTACT (9)
value PAN_LETT_OBLIQUE_FLATTENED (12)
value PAN_LETT_OBLIQUE_OFF_CENTER (14)
value PAN_LETT_OBLIQUE_ROUNDED (13)
value PAN_LETT_OBLIQUE_SQUARE (15)
value PAN_LETT_OBLIQUE_WEIGHTED (10)
value PAN_MIDLINE_CONSTANT_POINTED (9)
value PAN_MIDLINE_CONSTANT_SERIFED (10)
value PAN_MIDLINE_CONSTANT_TRIMMED (8)
value PAN_MIDLINE_HIGH_POINTED (6)
value PAN_MIDLINE_HIGH_SERIFED (7)
value PAN_MIDLINE_HIGH_TRIMMED (5)
value PAN_MIDLINE_INDEX (8)
value PAN_MIDLINE_LOW_POINTED (12)
value PAN_MIDLINE_LOW_SERIFED (13)
value PAN_MIDLINE_LOW_TRIMMED (11)
value PAN_MIDLINE_STANDARD_POINTED (3)
value PAN_MIDLINE_STANDARD_SERIFED (4)
value PAN_MIDLINE_STANDARD_TRIMMED (2)
value PAN_NO_FIT (1)
value PAN_PROPORTION_INDEX (3)
value PAN_PROP_CONDENSED (6)
value PAN_PROP_EVEN_WIDTH (4)
value PAN_PROP_EXPANDED (5)
value PAN_PROP_MODERN (3)
value PAN_PROP_MONOSPACED (9)
value PAN_PROP_OLD_STYLE (2)
value PAN_PROP_VERY_CONDENSED (8)
value PAN_PROP_VERY_EXPANDED (7)
value PAN_SERIFSTYLE_INDEX (1)
value PAN_SERIF_BONE (8)
value PAN_SERIF_COVE (2)
value PAN_SERIF_EXAGGERATED (9)
value PAN_SERIF_FLARED (14)
value PAN_SERIF_NORMAL_SANS (11)
value PAN_SERIF_OBTUSE_COVE (3)
value PAN_SERIF_OBTUSE_SANS (12)
value PAN_SERIF_OBTUSE_SQUARE_COVE (5)
value PAN_SERIF_PERP_SANS (13)
value PAN_SERIF_ROUNDED (15)
value PAN_SERIF_SQUARE (6)
value PAN_SERIF_SQUARE_COVE (4)
value PAN_SERIF_THIN (7)
value PAN_SERIF_TRIANGLE (10)
value PAN_STRAIGHT_ARMS_DOUBLE_SERIF (6)
value PAN_STRAIGHT_ARMS_HORZ (2)
value PAN_STRAIGHT_ARMS_SINGLE_SERIF (5)
value PAN_STRAIGHT_ARMS_VERT (4)
value PAN_STRAIGHT_ARMS_WEDGE (3)
value PAN_STROKEVARIATION_INDEX (5)
value PAN_STROKE_GRADUAL_DIAG (2)
value PAN_STROKE_GRADUAL_HORZ (5)
value PAN_STROKE_GRADUAL_TRAN (3)
value PAN_STROKE_GRADUAL_VERT (4)
value PAN_STROKE_INSTANT_VERT (8)
value PAN_STROKE_RAPID_HORZ (7)
value PAN_STROKE_RAPID_VERT (6)
value PAN_WEIGHT_BLACK (10)
value PAN_WEIGHT_BOLD (8)
value PAN_WEIGHT_BOOK (5)
value PAN_WEIGHT_DEMI (7)
value PAN_WEIGHT_HEAVY (9)
value PAN_WEIGHT_INDEX (2)
value PAN_WEIGHT_LIGHT (3)
value PAN_WEIGHT_MEDIUM (6)
value PAN_WEIGHT_NORD (11)
value PAN_WEIGHT_THIN (4)
value PAN_WEIGHT_VERY_LIGHT (2)
value PAN_XHEIGHT_CONSTANT_LARGE (4)
value PAN_XHEIGHT_CONSTANT_SMALL (2)
value PAN_XHEIGHT_CONSTANT_STD (3)
value PAN_XHEIGHT_DUCKING_LARGE (7)
value PAN_XHEIGHT_DUCKING_SMALL (5)
value PAN_XHEIGHT_DUCKING_STD (6)
value PAN_XHEIGHT_INDEX (9)
value PARAMFLAG_FHASCUSTDATA (( 0x40 ))
value PARAMFLAG_FHASDEFAULT (( 0x20 ))
value PARAMFLAG_FIN (( 0x1 ))
value PARAMFLAG_FLCID (( 0x4 ))
value PARAMFLAG_FOPT (( 0x10 ))
value PARAMFLAG_FOUT (( 0x2 ))
value PARAMFLAG_FRETVAL (( 0x8 ))
value PARAMFLAG_NONE (( 0 ))
value PARITY_EVEN (((WORD)0x0400))
value PARITY_MARK (((WORD)0x0800))
value PARITY_NONE (((WORD)0x0100))
value PARITY_ODD (((WORD)0x0200))
value PARITY_SPACE (((WORD)0x1000))
value PARKING_TOPOLOGY_POLICY_DISABLED (0)
value PARKING_TOPOLOGY_POLICY_ROUNDROBIN (1)
value PARKING_TOPOLOGY_POLICY_SEQUENTIAL (2)
value PARSE_DECODE (8)
value PARSE_ENCODE (7)
value PARTIITON_OS_DATA (0x29)
value PARTITION_BSP (0x2b)
value PARTITION_DM (0x54)
value PARTITION_DPP (0x2c)
value PARTITION_ENTRY_UNUSED (0x00)
value PARTITION_EXTENDED (0x05)
value PARTITION_EZDRIVE (0x55)
value PARTITION_GPT (0xEE)
value PARTITION_HUGE (0x06)
value PARTITION_IFS (0x07)
value PARTITION_LDM (0x42)
value PARTITION_MAIN_OS (0x28)
value PARTITION_MSFT_RECOVERY (0x27)
value PARTITION_NTFT (0x80)
value PARTITION_PREP (0x41)
value PARTITION_PRE_INSTALLED (0x2a)
value PARTITION_SPACES (0xE7)
value PARTITION_SPACES_DATA (0xD7)
value PARTITION_SYSTEM (0xEF)
value PARTITION_UNIX (0x63)
value PARTITION_WINDOWS_SYSTEM (0x2d)
value PASSEMBLY_DLL_REDIRECTION_DETAILED_INFORMATION (PASSEMBLY_FILE_DETAILED_INFORMATION)
value PASSIVE_LEVEL (0)
value PASSTHROUGH (19)
value PATCOPY ((DWORD)0x00F00021)
value PATINVERT ((DWORD)0x005A0049)
value PATPAINT ((DWORD)0x00FB0A09)
value PA_ACTIVATE (MA_ACTIVATE)
value PA_NOACTIVATE (MA_NOACTIVATE)
value PBTF_APMRESUMEFROMFAILURE (0x00000001)
value PBT_APMBATTERYLOW (0x0009)
value PBT_APMOEMEVENT (0x000B)
value PBT_APMPOWERSTATUSCHANGE (0x000A)
value PBT_APMQUERYSTANDBY (0x0001)
value PBT_APMQUERYSTANDBYFAILED (0x0003)
value PBT_APMQUERYSUSPEND (0x0000)
value PBT_APMQUERYSUSPENDFAILED (0x0002)
value PBT_APMRESUMEAUTOMATIC (0x0012)
value PBT_APMRESUMECRITICAL (0x0006)
value PBT_APMRESUMESTANDBY (0x0008)
value PBT_APMRESUMESUSPEND (0x0007)
value PBT_APMSTANDBY (0x0005)
value PBT_APMSUSPEND (0x0004)
value PBT_POWERSETTINGCHANGE (0x8013)
value PCASSEMBLY_DLL_REDIRECTION_DETAILED_INFORMATION (PCASSEMBLY_FILE_DETAILED_INFORMATION)
value PCF_DTRDSR (((DWORD)0x0001))
value PCF_INTTIMEOUTS (((DWORD)0x0080))
value PCF_PARITY_CHECK (((DWORD)0x0008))
value PCF_RLSD (((DWORD)0x0004))
value PCF_RTSCTS (((DWORD)0x0002))
value PCF_SETXCHAR (((DWORD)0x0020))
value PCF_SPECIALCHARS (((DWORD)0x0100))
value PCF_TOTALTIMEOUTS (((DWORD)0x0040))
value PCF_XONXOFF (((DWORD)0x0010))
value PCLEANUI ((SHTDN_REASON_FLAG_PLANNED | SHTDN_REASON_FLAG_CLEAN_UI))
value PC_EXPLICIT (0x02)
value PC_INTERIORS (128)
value PC_NOCOLLAPSE (0x04)
value PC_NONE (0)
value PC_PATHS (512)
value PC_POLYGON (1)
value PC_POLYPOLYGON (256)
value PC_RECTANGLE (2)
value PC_RESERVED (0x01)
value PC_SCANLINE (8)
value PC_STYLED (32)
value PC_TRAPEZOID (4)
value PC_WIDE (16)
value PC_WIDESTYLED (64)
value PC_WINDPOLYGON (4)
value PDCAP_WARM_EJECT_SUPPORTED (0x00000100)
value PDC_ARRIVAL (0x001)
value PDC_MAPPING_CHANGE (0x100)
value PDC_MODE_ASPECTRATIOPRESERVED (0x800)
value PDC_MODE_CENTERED (0x080)
value PDC_MODE_DEFAULT (0x040)
value PDC_ORIGIN (0x400)
value PDC_REMOVAL (0x002)
value PDC_RESOLUTION (0x200)
value PDERR_CREATEICFAILURE (0x100A)
value PDERR_DEFAULTDIFFERENT (0x100C)
value PDERR_DNDMMISMATCH (0x1009)
value PDERR_GETDEVMODEFAIL (0x1005)
value PDERR_INITFAILURE (0x1006)
value PDERR_LOADDRVFAILURE (0x1004)
value PDERR_NODEFAULTPRN (0x1008)
value PDERR_NODEVICES (0x1007)
value PDERR_PARSEFAILURE (0x1002)
value PDERR_PRINTERCODES (0x1000)
value PDERR_PRINTERNOTFOUND (0x100B)
value PDERR_RETDEFFAILURE (0x1003)
value PDERR_SETUPFAILURE (0x1001)
value PDEVICESIZE (26)
value PDIRTYUI ((SHTDN_REASON_FLAG_PLANNED | SHTDN_REASON_FLAG_DIRTY_UI))
value PD_ALLPAGES (0x00000000)
value PD_COLLATE (0x00000010)
value PD_CURRENTPAGE (0x00400000)
value PD_DISABLEPRINTTOFILE (0x00080000)
value PD_ENABLEPRINTHOOK (0x00001000)
value PD_ENABLEPRINTTEMPLATE (0x00004000)
value PD_ENABLEPRINTTEMPLATEHANDLE (0x00010000)
value PD_ENABLESETUPHOOK (0x00002000)
value PD_ENABLESETUPTEMPLATE (0x00008000)
value PD_ENABLESETUPTEMPLATEHANDLE (0x00020000)
value PD_EXCLUSIONFLAGS (0x01000000)
value PD_EXCL_COPIESANDCOLLATE ((DM_COPIES | DM_COLLATE))
value PD_HIDEPRINTTOFILE (0x00100000)
value PD_NOCURRENTPAGE (0x00800000)
value PD_NONETWORKBUTTON (0x00200000)
value PD_NOPAGENUMS (0x00000008)
value PD_NOSELECTION (0x00000004)
value PD_NOWARNING (0x00000080)
value PD_PAGENUMS (0x00000002)
value PD_PRINTSETUP (0x00000040)
value PD_PRINTTOFILE (0x00000020)
value PD_RESULT_APPLY (2)
value PD_RESULT_CANCEL (0)
value PD_RESULT_PRINT (1)
value PD_RETURNDC (0x00000100)
value PD_RETURNDEFAULT (0x00000400)
value PD_RETURNIC (0x00000200)
value PD_SELECTION (0x00000001)
value PD_SHOWHELP (0x00000800)
value PD_USEDEVMODECOPIES (0x00040000)
value PD_USEDEVMODECOPIESANDCOLLATE (0x00040000)
value PD_USELARGETEMPLATE (0x10000000)
value PEERDIST_ERROR_ALREADY_COMPLETED (4060)
value PEERDIST_ERROR_ALREADY_EXISTS (4058)
value PEERDIST_ERROR_ALREADY_INITIALIZED (4055)
value PEERDIST_ERROR_CANNOT_PARSE_CONTENTINFO (4051)
value PEERDIST_ERROR_CONTENTINFO_VERSION_UNSUPPORTED (4050)
value PEERDIST_ERROR_INVALIDATED (4057)
value PEERDIST_ERROR_INVALID_CONFIGURATION (4063)
value PEERDIST_ERROR_MISSING_DATA (4052)
value PEERDIST_ERROR_NOT_INITIALIZED (4054)
value PEERDIST_ERROR_NOT_LICENSED (4064)
value PEERDIST_ERROR_NO_MORE (4053)
value PEERDIST_ERROR_OPERATION_NOTFOUND (4059)
value PEERDIST_ERROR_OUT_OF_BOUNDS (4061)
value PEERDIST_ERROR_SERVICE_UNAVAILABLE (4065)
value PEERDIST_ERROR_SHUTDOWN_IN_PROGRESS (4056)
value PEERDIST_ERROR_TRUST_FAILURE (4066)
value PEERDIST_ERROR_VERSION_UNSUPPORTED (4062)
value PEER_E_ALREADY_LISTENING (_HRESULT_TYPEDEF_(0x80630107L))
value PEER_E_CANNOT_CONVERT_PEER_NAME (_HRESULT_TYPEDEF_(0x80634001L))
value PEER_E_CANNOT_START_SERVICE (_HRESULT_TYPEDEF_(0x80630003L))
value PEER_E_CERT_STORE_CORRUPTED (_HRESULT_TYPEDEF_(0x80630801L))
value PEER_E_CHAIN_TOO_LONG (_HRESULT_TYPEDEF_(0x80630703L))
value PEER_E_CIRCULAR_CHAIN_DETECTED (_HRESULT_TYPEDEF_(0x80630706L))
value PEER_E_CLASSIFIER_TOO_LONG (_HRESULT_TYPEDEF_(0x80630201L))
value PEER_E_CLOUD_NAME_AMBIGUOUS (_HRESULT_TYPEDEF_(0x80631005L))
value PEER_E_CONNECTION_FAILED (_HRESULT_TYPEDEF_(0x80630109L))
value PEER_E_CONNECTION_NOT_AUTHENTICATED (_HRESULT_TYPEDEF_(0x8063010AL))
value PEER_E_CONNECTION_NOT_FOUND (_HRESULT_TYPEDEF_(0x80630103L))
value PEER_E_CONNECTION_REFUSED (_HRESULT_TYPEDEF_(0x8063010BL))
value PEER_E_CONNECT_SELF (_HRESULT_TYPEDEF_(0x80630106L))
value PEER_E_CONTACT_NOT_FOUND (_HRESULT_TYPEDEF_(0x80636001L))
value PEER_E_DATABASE_ACCESSDENIED (_HRESULT_TYPEDEF_(0x80630302L))
value PEER_E_DATABASE_ALREADY_PRESENT (_HRESULT_TYPEDEF_(0x80630305L))
value PEER_E_DATABASE_NOT_PRESENT (_HRESULT_TYPEDEF_(0x80630306L))
value PEER_E_DBINITIALIZATION_FAILED (_HRESULT_TYPEDEF_(0x80630303L))
value PEER_E_DBNAME_CHANGED (_HRESULT_TYPEDEF_(0x80630011L))
value PEER_E_DEFERRED_VALIDATION (_HRESULT_TYPEDEF_(0x80632030L))
value PEER_E_DUPLICATE_GRAPH (_HRESULT_TYPEDEF_(0x80630012L))
value PEER_E_EVENT_HANDLE_NOT_FOUND (_HRESULT_TYPEDEF_(0x80630501L))
value PEER_E_FW_BLOCKED_BY_POLICY (_HRESULT_TYPEDEF_(0x80637009L))
value PEER_E_FW_BLOCKED_BY_SHIELDS_UP (_HRESULT_TYPEDEF_(0x8063700AL))
value PEER_E_FW_DECLINED (_HRESULT_TYPEDEF_(0x8063700BL))
value PEER_E_FW_EXCEPTION_DISABLED (_HRESULT_TYPEDEF_(0x80637008L))
value PEER_E_GRAPH_IN_USE (_HRESULT_TYPEDEF_(0x80630015L))
value PEER_E_GRAPH_NOT_READY (_HRESULT_TYPEDEF_(0x80630013L))
value PEER_E_GRAPH_SHUTTING_DOWN (_HRESULT_TYPEDEF_(0x80630014L))
value PEER_E_GROUPS_EXIST (_HRESULT_TYPEDEF_(0x80630204L))
value PEER_E_GROUP_IN_USE (_HRESULT_TYPEDEF_(0x80632092L))
value PEER_E_GROUP_NOT_READY (_HRESULT_TYPEDEF_(0x80632091L))
value PEER_E_IDENTITY_DELETED (_HRESULT_TYPEDEF_(0x806320A0L))
value PEER_E_IDENTITY_NOT_FOUND (_HRESULT_TYPEDEF_(0x80630401L))
value PEER_E_INVALID_ADDRESS (_HRESULT_TYPEDEF_(0x80637007L))
value PEER_E_INVALID_ATTRIBUTES (_HRESULT_TYPEDEF_(0x80630602L))
value PEER_E_INVALID_CLASSIFIER (_HRESULT_TYPEDEF_(0x80632060L))
value PEER_E_INVALID_CLASSIFIER_PROPERTY (_HRESULT_TYPEDEF_(0x80632072L))
value PEER_E_INVALID_CREDENTIAL (_HRESULT_TYPEDEF_(0x80632082L))
value PEER_E_INVALID_CREDENTIAL_INFO (_HRESULT_TYPEDEF_(0x80632081L))
value PEER_E_INVALID_DATABASE (_HRESULT_TYPEDEF_(0x80630016L))
value PEER_E_INVALID_FRIENDLY_NAME (_HRESULT_TYPEDEF_(0x80632070L))
value PEER_E_INVALID_GRAPH (_HRESULT_TYPEDEF_(0x80630010L))
value PEER_E_INVALID_GROUP (_HRESULT_TYPEDEF_(0x80632093L))
value PEER_E_INVALID_GROUP_PROPERTIES (_HRESULT_TYPEDEF_(0x80632040L))
value PEER_E_INVALID_PEER_HOST_NAME (_HRESULT_TYPEDEF_(0x80634002L))
value PEER_E_INVALID_PEER_NAME (_HRESULT_TYPEDEF_(0x80632050L))
value PEER_E_INVALID_RECORD (_HRESULT_TYPEDEF_(0x80632010L))
value PEER_E_INVALID_RECORD_EXPIRATION (_HRESULT_TYPEDEF_(0x80632080L))
value PEER_E_INVALID_RECORD_SIZE (_HRESULT_TYPEDEF_(0x80632083L))
value PEER_E_INVALID_ROLE_PROPERTY (_HRESULT_TYPEDEF_(0x80632071L))
value PEER_E_INVALID_SEARCH (_HRESULT_TYPEDEF_(0x80630601L))
value PEER_E_INVALID_TIME_PERIOD (_HRESULT_TYPEDEF_(0x80630705L))
value PEER_E_INVITATION_NOT_TRUSTED (_HRESULT_TYPEDEF_(0x80630701L))
value PEER_E_INVITE_CANCELLED (_HRESULT_TYPEDEF_(0x80637000L))
value PEER_E_INVITE_RESPONSE_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x80637001L))
value PEER_E_MAX_RECORD_SIZE_EXCEEDED (_HRESULT_TYPEDEF_(0x80630304L))
value PEER_E_NODE_NOT_FOUND (_HRESULT_TYPEDEF_(0x80630108L))
value PEER_E_NOT_AUTHORIZED (_HRESULT_TYPEDEF_(0x80632020L))
value PEER_E_NOT_INITIALIZED (_HRESULT_TYPEDEF_(0x80630002L))
value PEER_E_NOT_LICENSED (_HRESULT_TYPEDEF_(0x80630004L))
value PEER_E_NOT_SIGNED_IN (_HRESULT_TYPEDEF_(0x80637003L))
value PEER_E_NO_CLOUD (_HRESULT_TYPEDEF_(0x80631001L))
value PEER_E_NO_KEY_ACCESS (_HRESULT_TYPEDEF_(0x80630203L))
value PEER_E_NO_MEMBERS_FOUND (_HRESULT_TYPEDEF_(0x80632094L))
value PEER_E_NO_MEMBER_CONNECTIONS (_HRESULT_TYPEDEF_(0x80632095L))
value PEER_E_NO_MORE (_HRESULT_TYPEDEF_(0x80634003L))
value PEER_E_PASSWORD_DOES_NOT_MEET_POLICY (_HRESULT_TYPEDEF_(0x80632021L))
value PEER_E_PNRP_DUPLICATE_PEER_NAME (_HRESULT_TYPEDEF_(0x80634005L))
value PEER_E_PRIVACY_DECLINED (_HRESULT_TYPEDEF_(0x80637004L))
value PEER_E_RECORD_NOT_FOUND (_HRESULT_TYPEDEF_(0x80630301L))
value PEER_E_SERVICE_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x806320A1L))
value PEER_E_TIMEOUT (_HRESULT_TYPEDEF_(0x80637005L))
value PEER_E_TOO_MANY_ATTRIBUTES (_HRESULT_TYPEDEF_(0x80630017L))
value PEER_E_TOO_MANY_IDENTITIES (_HRESULT_TYPEDEF_(0x80630202L))
value PEER_E_UNABLE_TO_LISTEN (_HRESULT_TYPEDEF_(0x80632096L))
value PEER_E_UNSUPPORTED_VERSION (_HRESULT_TYPEDEF_(0x80632090L))
value PEER_S_ALREADY_A_MEMBER (_HRESULT_TYPEDEF_(0x00630006L))
value PEER_S_ALREADY_CONNECTED (_HRESULT_TYPEDEF_(0x00632000L))
value PEER_S_GRAPH_DATA_CREATED (_HRESULT_TYPEDEF_(0x00630001L))
value PEER_S_NO_CONNECTIVITY (_HRESULT_TYPEDEF_(0x00630005L))
value PEER_S_NO_EVENT_DATA (_HRESULT_TYPEDEF_(0x00630002L))
value PEER_S_SUBSCRIPTION_EXISTS (_HRESULT_TYPEDEF_(0x00636000L))
value PENARBITRATIONTYPE_FIS (0x0002)
value PENARBITRATIONTYPE_MAX (0x0004)
value PENARBITRATIONTYPE_NONE (0x0000)
value PENARBITRATIONTYPE_SPT (0x0003)
value PENVISUALIZATION_CURSOR (0x0020)
value PENVISUALIZATION_DOUBLETAP (0x0002)
value PENVISUALIZATION_OFF (0x0000)
value PENVISUALIZATION_ON (0x0023)
value PENVISUALIZATION_TAP (0x0001)
value PEN_FLAG_BARREL (0x00000001)
value PEN_FLAG_ERASER (0x00000004)
value PEN_FLAG_INVERTED (0x00000002)
value PEN_FLAG_NONE (0x00000000)
value PEN_MASK_NONE (0x00000000)
value PEN_MASK_PRESSURE (0x00000001)
value PEN_MASK_ROTATION (0x00000002)
value PEN_MASK_TILT_X (0x00000004)
value PEN_MASK_TILT_Y (0x00000008)
value PERFORMANCE_DATA_VERSION (1)
value PERFSTATE_POLICY_CHANGE_DECREASE_MAX (PERFSTATE_POLICY_CHANGE_ROCKET)
value PERFSTATE_POLICY_CHANGE_IDEAL (0)
value PERFSTATE_POLICY_CHANGE_IDEAL_AGGRESSIVE (3)
value PERFSTATE_POLICY_CHANGE_INCREASE_MAX (PERFSTATE_POLICY_CHANGE_IDEAL_AGGRESSIVE)
value PERFSTATE_POLICY_CHANGE_ROCKET (2)
value PERFSTATE_POLICY_CHANGE_SINGLE (1)
value PERF_AVERAGE_BASE ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_BASE | PERF_DISPLAY_NOSHOW | 0x00000002))
value PERF_AVERAGE_BULK ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_FRACTION | PERF_DISPLAY_NOSHOW))
value PERF_AVERAGE_TIMER ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_FRACTION | PERF_DISPLAY_SECONDS))
value PERF_COUNTER_BASE (0x00030000)
value PERF_COUNTER_BULK_COUNT ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_RATE | PERF_TIMER_TICK | PERF_DELTA_COUNTER | PERF_DISPLAY_PER_SEC))
value PERF_COUNTER_COUNTER ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_RATE | PERF_TIMER_TICK | PERF_DELTA_COUNTER | PERF_DISPLAY_PER_SEC))
value PERF_COUNTER_DELTA ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_VALUE | PERF_DELTA_COUNTER | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_ELAPSED (0x00040000)
value PERF_COUNTER_FRACTION (0x00020000)
value PERF_COUNTER_HISTOGRAM (0x00060000)
value PERF_COUNTER_HISTOGRAM_TYPE (0x80000000)
value PERF_COUNTER_LARGE_DELTA ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_VALUE | PERF_DELTA_COUNTER | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_LARGE_QUEUELEN_TYPE ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_QUEUELEN | PERF_TIMER_TICK | PERF_DELTA_COUNTER | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_LARGE_RAWCOUNT ((PERF_SIZE_LARGE | PERF_TYPE_NUMBER | PERF_NUMBER_DECIMAL | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_LARGE_RAWCOUNT_HEX ((PERF_SIZE_LARGE | PERF_TYPE_NUMBER | PERF_NUMBER_HEX | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_MULTI_BASE ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_BASE | PERF_MULTI_COUNTER | PERF_DISPLAY_NOSHOW))
value PERF_COUNTER_MULTI_TIMER ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_RATE | PERF_DELTA_COUNTER | PERF_TIMER_TICK | PERF_MULTI_COUNTER | PERF_DISPLAY_PERCENT))
value PERF_COUNTER_MULTI_TIMER_INV ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_RATE | PERF_DELTA_COUNTER | PERF_MULTI_COUNTER | PERF_TIMER_TICK | PERF_INVERSE_COUNTER | PERF_DISPLAY_PERCENT))
value PERF_COUNTER_NODATA ((PERF_SIZE_ZERO | PERF_DISPLAY_NOSHOW))
value PERF_COUNTER_OBJ_TIME_QUEUELEN_TYPE ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_QUEUELEN | PERF_OBJECT_TIMER | PERF_DELTA_COUNTER | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_PRECISION (0x00070000)
value PERF_COUNTER_QUEUELEN (0x00050000)
value PERF_COUNTER_QUEUELEN_TYPE ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_QUEUELEN | PERF_TIMER_TICK | PERF_DELTA_COUNTER | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_RATE (0x00010000)
value PERF_COUNTER_RAWCOUNT ((PERF_SIZE_DWORD | PERF_TYPE_NUMBER | PERF_NUMBER_DECIMAL | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_RAWCOUNT_HEX ((PERF_SIZE_DWORD | PERF_TYPE_NUMBER | PERF_NUMBER_HEX | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_TEXT ((PERF_SIZE_VARIABLE_LEN | PERF_TYPE_TEXT | PERF_TEXT_UNICODE | PERF_DISPLAY_NO_SUFFIX))
value PERF_COUNTER_TIMER ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_RATE | PERF_TIMER_TICK | PERF_DELTA_COUNTER | PERF_DISPLAY_PERCENT))
value PERF_COUNTER_TIMER_INV ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_RATE | PERF_TIMER_TICK | PERF_DELTA_COUNTER | PERF_INVERSE_COUNTER | PERF_DISPLAY_PERCENT))
value PERF_COUNTER_VALUE (0x00000000)
value PERF_DATA_REVISION (1)
value PERF_DATA_VERSION (1)
value PERF_DELTA_BASE (0x00800000)
value PERF_DELTA_COUNTER (0x00400000)
value PERF_DETAIL_ADVANCED (200)
value PERF_DETAIL_EXPERT (300)
value PERF_DETAIL_NOVICE (100)
value PERF_DETAIL_WIZARD (400)
value PERF_DISPLAY_NOSHOW (0x40000000)
value PERF_DISPLAY_NO_SUFFIX (0x00000000)
value PERF_DISPLAY_PERCENT (0x20000000)
value PERF_DISPLAY_PER_SEC (0x10000000)
value PERF_DISPLAY_SECONDS (0x30000000)
value PERF_ELAPSED_TIME ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_ELAPSED | PERF_OBJECT_TIMER | PERF_DISPLAY_SECONDS))
value PERF_INVERSE_COUNTER (0x01000000)
value PERF_LARGE_RAW_BASE ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_BASE | PERF_DISPLAY_NOSHOW ))
value PERF_LARGE_RAW_FRACTION ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_FRACTION | PERF_DISPLAY_PERCENT))
value PERF_METADATA_MULTIPLE_INSTANCES ((-2))
value PERF_METADATA_NO_INSTANCES ((-3))
value PERF_MULTI_COUNTER (0x02000000)
value PERF_NO_INSTANCES ((-1))
value PERF_NO_UNIQUE_ID (-1)
value PERF_NUMBER_DECIMAL (0x00010000)
value PERF_NUMBER_HEX (0x00000000)
value PERF_OBJECT_TIMER (0x00200000)
value PERF_OBJ_TIME_TIMER ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_RATE | PERF_OBJECT_TIMER | PERF_DELTA_COUNTER | PERF_DISPLAY_PERCENT))
value PERF_PRECISION_OBJECT_TIMER ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_PRECISION | PERF_OBJECT_TIMER | PERF_DELTA_COUNTER | PERF_DISPLAY_PERCENT ))
value PERF_PRECISION_SYSTEM_TIMER ((PERF_SIZE_LARGE | PERF_TYPE_COUNTER | PERF_COUNTER_PRECISION | PERF_TIMER_TICK | PERF_DELTA_COUNTER | PERF_DISPLAY_PERCENT ))
value PERF_PRECISION_TIMESTAMP (PERF_LARGE_RAW_BASE)
value PERF_RAW_BASE ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_BASE | PERF_DISPLAY_NOSHOW | 0x00000003))
value PERF_RAW_FRACTION ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_FRACTION | PERF_DISPLAY_PERCENT))
value PERF_SAMPLE_BASE ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_BASE | PERF_DISPLAY_NOSHOW | 0x00000001))
value PERF_SAMPLE_COUNTER ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_RATE | PERF_TIMER_TICK | PERF_DELTA_COUNTER | PERF_DISPLAY_NO_SUFFIX))
value PERF_SAMPLE_FRACTION ((PERF_SIZE_DWORD | PERF_TYPE_COUNTER | PERF_COUNTER_FRACTION | PERF_DELTA_COUNTER | PERF_DELTA_BASE | PERF_DISPLAY_PERCENT))
value PERF_SIZE_DWORD (0x00000000)
value PERF_SIZE_LARGE (0x00000100)
value PERF_SIZE_VARIABLE_LEN (0x00000300)
value PERF_SIZE_ZERO (0x00000200)
value PERF_TEXT_ASCII (0x00010000)
value PERF_TEXT_UNICODE (0x00000000)
value PERF_TIMER_TICK (0x00000000)
value PERF_TYPE_COUNTER (0x00000400)
value PERF_TYPE_NUMBER (0x00000000)
value PERF_TYPE_TEXT (0x00000800)
value PERF_TYPE_ZERO (0x00000C00)
value PERSISTENT_VOLUME_STATE_BACKED_BY_WIM ((0x00000040))
value PERSISTENT_VOLUME_STATE_CHKDSK_RAN_ONCE ((0x00000400))
value PERSISTENT_VOLUME_STATE_CONTAINS_BACKING_WIM ((0x00000020))
value PERSISTENT_VOLUME_STATE_DAX_FORMATTED ((0x00001000))
value PERSISTENT_VOLUME_STATE_GLOBAL_METADATA_NO_SEEK_PENALTY ((0x00000004))
value PERSISTENT_VOLUME_STATE_LOCAL_METADATA_NO_SEEK_PENALTY ((0x00000008))
value PERSISTENT_VOLUME_STATE_MODIFIED_BY_CHKDSK ((0x00000800))
value PERSISTENT_VOLUME_STATE_NO_HEAT_GATHERING ((0x00000010))
value PERSISTENT_VOLUME_STATE_NO_WRITE_AUTO_TIERING ((0x00000080))
value PERSISTENT_VOLUME_STATE_REALLOCATE_ALL_DATA_WRITES ((0x00000200))
value PERSISTENT_VOLUME_STATE_SHORT_NAME_CREATION_DISABLED ((0x00000001))
value PERSISTENT_VOLUME_STATE_TXF_DISABLED ((0x00000100))
value PERSISTENT_VOLUME_STATE_VOLUME_SCRUB_DISABLED ((0x00000002))
value PERSIST_E_NOTSELFSIZING (_HRESULT_TYPEDEF_(0x800B000BL))
value PERSIST_E_SIZEDEFINITE (_HRESULT_TYPEDEF_(0x800B0009L))
value PERSIST_E_SIZEINDEFINITE (_HRESULT_TYPEDEF_(0x800B000AL))
value PFD_DEPTH_DONTCARE (0x20000000)
value PFD_DOUBLEBUFFER (0x00000001)
value PFD_DOUBLEBUFFER_DONTCARE (0x40000000)
value PFD_DRAW_TO_BITMAP (0x00000008)
value PFD_DRAW_TO_WINDOW (0x00000004)
value PFD_GENERIC_ACCELERATED (0x00001000)
value PFD_GENERIC_FORMAT (0x00000040)
value PFD_MAIN_PLANE (0)
value PFD_NEED_PALETTE (0x00000080)
value PFD_NEED_SYSTEM_PALETTE (0x00000100)
value PFD_OVERLAY_PLANE (1)
value PFD_STEREO (0x00000002)
value PFD_STEREO_DONTCARE (0x80000000)
value PFD_SUPPORT_COMPOSITION (0x00008000)
value PFD_SUPPORT_DIRECTDRAW (0x00002000)
value PFD_SUPPORT_GDI (0x00000010)
value PFD_SUPPORT_OPENGL (0x00000020)
value PFD_SWAP_COPY (0x00000400)
value PFD_SWAP_EXCHANGE (0x00000200)
value PFD_SWAP_LAYER_BUFFERS (0x00000800)
value PFD_TYPE_COLORINDEX (1)
value PFD_TYPE_RGBA (0)
value PFD_UNDERLAY_PLANE ((-1))
value PFL_HIDDEN (0x00000004)
value PFL_MATCHES_PROTOCOL_ZERO (0x00000008)
value PFL_MULTIPLE_PROTO_ENTRIES (0x00000001)
value PFL_NETWORKDIRECT_PROVIDER (0x00000010)
value PFL_RECOMMENDED_PROTO_ENTRY (0x00000002)
value PFORCEINLINE (FORCEINLINE)
value PF_ALPHA_BYTE_INSTRUCTIONS (5)
value PF_APPLETALK (AF_APPLETALK)
value PF_ARM_DIVIDE_INSTRUCTION_AVAILABLE (24)
value PF_ARM_EXTERNAL_CACHE_AVAILABLE (26)
value PF_ARM_FMAC_INSTRUCTIONS_AVAILABLE (27)
value PF_ARM_NEON_INSTRUCTIONS_AVAILABLE (19)
value PF_ATM (AF_ATM)
value PF_AVX_INSTRUCTIONS_AVAILABLE (39)
value PF_BAN (AF_BAN)
value PF_BTH (AF_BTH)
value PF_CCITT (AF_CCITT)
value PF_CHANNELS_ENABLED (16)
value PF_CHAOS (AF_CHAOS)
value PF_COMPARE_EXCHANGE_DOUBLE (2)
value PF_DATAKIT (AF_DATAKIT)
value PF_DLI (AF_DLI)
value PF_ECMA (AF_ECMA)
value PF_ERMS_AVAILABLE (42)
value PF_FASTFAIL_AVAILABLE (23)
value PF_FIREFOX (AF_FIREFOX)
value PF_FLOATING_POINT_EMULATED (1)
value PF_FLOATING_POINT_PRECISION_ERRATA (0)
value PF_HYLINK (AF_HYLINK)
value PF_IMPLINK (AF_IMPLINK)
value PF_INET (AF_INET)
value PF_IPX (AF_IPX)
value PF_ISO (AF_ISO)
value PF_LAT (AF_LAT)
value PF_MAX (AF_MAX)
value PF_MMX_INSTRUCTIONS_AVAILABLE (3)
value PF_MONITORX_INSTRUCTION_AVAILABLE (35)
value PF_NON_TEMPORAL_LEVEL_ALL (_MM_HINT_NTA)
value PF_NS (AF_NS)
value PF_NX_ENABLED (12)
value PF_OSI (AF_OSI)
value PF_PAE_ENABLED (9)
value PF_PUP (AF_PUP)
value PF_RDPID_INSTRUCTION_AVAILABLE (33)
value PF_RDRAND_INSTRUCTION_AVAILABLE (28)
value PF_RDTSCP_INSTRUCTION_AVAILABLE (32)
value PF_RDTSC_INSTRUCTION_AVAILABLE (8)
value PF_RDWRFSGSBASE_AVAILABLE (22)
value PF_SECOND_LEVEL_ADDRESS_TRANSLATION (20)
value PF_SNA (AF_SNA)
value PF_SSE_DAZ_MODE_AVAILABLE (11)
value PF_UNIX (AF_UNIX)
value PF_UNSPEC (AF_UNSPEC)
value PF_VIRT_FIRMWARE_ENABLED (21)
value PF_VOICEVIEW (AF_VOICEVIEW)
value PF_XMMI_INSTRUCTIONS_AVAILABLE (6)
value PF_XSAVE_ENABLED (17)
value PGET_MODULE_HANDLE_EX (PGET_MODULE_HANDLE_EXA)
value PHYSICALHEIGHT (111)
value PHYSICALOFFSETX (112)
value PHYSICALOFFSETY (113)
value PHYSICALWIDTH (110)
value PIDDI_THUMBNAIL (0x00000002L)
value PIDDSI_BYTECOUNT (0x00000004)
value PIDDSI_CATEGORY (0x00000002)
value PIDDSI_COMPANY (0x0000000F)
value PIDDSI_DOCPARTS (0x0000000D)
value PIDDSI_HEADINGPAIR (0x0000000C)
value PIDDSI_HIDDENCOUNT (0x00000009)
value PIDDSI_LINECOUNT (0x00000005)
value PIDDSI_LINKSDIRTY (0x00000010)
value PIDDSI_MANAGER (0x0000000E)
value PIDDSI_MMCLIPCOUNT (0x0000000A)
value PIDDSI_NOTECOUNT (0x00000008)
value PIDDSI_PARCOUNT (0x00000006)
value PIDDSI_PRESFORMAT (0x00000003)
value PIDDSI_SCALE (0x0000000B)
value PIDDSI_SLIDECOUNT (0x00000007)
value PIDMSI_COPYRIGHT (0x0000000BL)
value PIDMSI_EDITOR (0x00000002L)
value PIDMSI_OWNER (0x00000008L)
value PIDMSI_PRODUCTION (0x0000000AL)
value PIDMSI_PROJECT (0x00000006L)
value PIDMSI_RATING (0x00000009L)
value PIDMSI_SEQUENCE_NO (0x00000005L)
value PIDMSI_SOURCE (0x00000004L)
value PIDMSI_STATUS (0x00000007L)
value PIDMSI_SUPPLIER (0x00000003L)
value PIDSI_APPNAME (0x00000012L)
value PIDSI_AUTHOR (0x00000004L)
value PIDSI_CHARCOUNT (0x00000010L)
value PIDSI_COMMENTS (0x00000006L)
value PIDSI_DOC_SECURITY (0x00000013L)
value PIDSI_KEYWORDS (0x00000005L)
value PIDSI_LASTAUTHOR (0x00000008L)
value PIDSI_REVNUMBER (0x00000009L)
value PIDSI_SUBJECT (0x00000003L)
value PIDSI_TEMPLATE (0x00000007L)
value PIDSI_THUMBNAIL (0x00000011L)
value PIDSI_TITLE (0x00000002L)
value PID_BEHAVIOR (( 0x80000003 ))
value PID_CODEPAGE (( 0x1 ))
value PID_DICTIONARY (( 0 ))
value PID_FIRST_USABLE (( 0x2 ))
value PID_LOCALE (( 0x80000000 ))
value PID_MIN_READONLY (( 0x80000000 ))
value PID_MODIFY_TIME (( 0x80000001 ))
value PID_SECURITY (( 0x80000002 ))
value PIPE_ACCEPT_REMOTE_CLIENTS (0x00000000)
value PIPE_ACCESS_DUPLEX (0x00000003)
value PIPE_ACCESS_INBOUND (0x00000001)
value PIPE_ACCESS_OUTBOUND (0x00000002)
value PIPE_CLIENT_END (0x00000000)
value PIPE_NOWAIT (0x00000001)
value PIPE_READMODE_BYTE (0x00000000)
value PIPE_READMODE_MESSAGE (0x00000002)
value PIPE_REJECT_REMOTE_CLIENTS (0x00000008)
value PIPE_SERVER_END (0x00000001)
value PIPE_TYPE_BYTE (0x00000000)
value PIPE_TYPE_MESSAGE (0x00000004)
value PIPE_UNLIMITED_INSTANCES (255)
value PIPE_WAIT (0x00000000)
value PI_DOCFILECLSIDLOOKUP (32)
value PKCS_ATTRIBUTE (((LPCSTR) 22))
value PKCS_ATTRIBUTES (((LPCSTR) 48))
value PKCS_CONTENT_INFO (((LPCSTR) 33))
value PKCS_CONTENT_INFO_SEQUENCE_OF_ANY (((LPCSTR) 23))
value PKCS_CTL (((LPCSTR) 37))
value PKCS_ENCRYPTED_PRIVATE_KEY_INFO (((LPCSTR) 45))
value PKCS_PRIVATE_KEY_INFO (((LPCSTR) 44))
value PKCS_RSAES_OAEP_PARAMETERS (((LPCSTR) 76))
value PKCS_RSA_PRIVATE_KEY (((LPCSTR) 43))
value PKCS_RSA_SSA_PSS_PARAMETERS (((LPCSTR) 75))
value PKCS_RSA_SSA_PSS_TRAILER_FIELD_BC (1)
value PKCS_SMIME_CAPABILITIES (((LPCSTR) 42))
value PKCS_SORTED_CTL (((LPCSTR) 49))
value PKCS_TIME_REQUEST (((LPCSTR) 18))
value PKCS_UTC_TIME (((LPCSTR) 17))
value PLAINTEXTKEYBLOB (0x8)
value PLANES (14)
value PLA_E_CABAPI_FAILURE (_HRESULT_TYPEDEF_(0x80300113L))
value PLA_E_CONFLICT_INCL_EXCL_API (_HRESULT_TYPEDEF_(0x80300105L))
value PLA_E_CREDENTIALS_REQUIRED (_HRESULT_TYPEDEF_(0x80300103L))
value PLA_E_DCS_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x803000B7L))
value PLA_E_DCS_IN_USE (_HRESULT_TYPEDEF_(0x803000AAL))
value PLA_E_DCS_NOT_FOUND (_HRESULT_TYPEDEF_(0x80300002L))
value PLA_E_DCS_NOT_RUNNING (_HRESULT_TYPEDEF_(0x80300104L))
value PLA_E_DCS_SINGLETON_REQUIRED (_HRESULT_TYPEDEF_(0x80300102L))
value PLA_E_DCS_START_WAIT_TIMEOUT (_HRESULT_TYPEDEF_(0x8030010AL))
value PLA_E_DC_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x80300109L))
value PLA_E_DC_START_WAIT_TIMEOUT (_HRESULT_TYPEDEF_(0x8030010BL))
value PLA_E_EXE_ALREADY_CONFIGURED (_HRESULT_TYPEDEF_(0x80300107L))
value PLA_E_EXE_FULL_PATH_REQUIRED (_HRESULT_TYPEDEF_(0x8030010EL))
value PLA_E_EXE_PATH_NOT_VALID (_HRESULT_TYPEDEF_(0x80300108L))
value PLA_E_INVALID_SESSION_NAME (_HRESULT_TYPEDEF_(0x8030010FL))
value PLA_E_NETWORK_EXE_NOT_VALID (_HRESULT_TYPEDEF_(0x80300106L))
value PLA_E_NO_DUPLICATES (_HRESULT_TYPEDEF_(0x8030010DL))
value PLA_E_NO_MIN_DISK (_HRESULT_TYPEDEF_(0x80300070L))
value PLA_E_PLA_CHANNEL_NOT_ENABLED (_HRESULT_TYPEDEF_(0x80300110L))
value PLA_E_PROPERTY_CONFLICT (_HRESULT_TYPEDEF_(0x80300101L))
value PLA_E_REPORT_WAIT_TIMEOUT (_HRESULT_TYPEDEF_(0x8030010CL))
value PLA_E_RULES_MANAGER_FAILED (_HRESULT_TYPEDEF_(0x80300112L))
value PLA_E_TASKSCHED_CHANNEL_NOT_ENABLED (_HRESULT_TYPEDEF_(0x80300111L))
value PLA_E_TOO_MANY_FOLDERS (_HRESULT_TYPEDEF_(0x80300045L))
value PLA_S_PROPERTY_IGNORED (_HRESULT_TYPEDEF_(0x00300100L))
value PMB_ACTIVE (0x00000001)
value PME_CURRENT_VERSION (1)
value PME_FAILFAST_ON_COMMIT_FAIL_DISABLE (0x0)
value PME_FAILFAST_ON_COMMIT_FAIL_ENABLE (0x1)
value PM_NOREMOVE (0x0000)
value PM_NOYIELD (0x0002)
value PM_REMOVE (0x0001)
value POINTER_DEVICE_PRODUCT_STRING_MAX (520)
value POINTER_FLAG_CANCELED (0x00008000)
value POINTER_FLAG_CAPTURECHANGED (0x00200000)
value POINTER_FLAG_CONFIDENCE (0x00004000)
value POINTER_FLAG_DOWN (0x00010000)
value POINTER_FLAG_FIFTHBUTTON (0x00000100)
value POINTER_FLAG_FIRSTBUTTON (0x00000010)
value POINTER_FLAG_FOURTHBUTTON (0x00000080)
value POINTER_FLAG_HASTRANSFORM (0x00400000)
value POINTER_FLAG_HWHEEL (0x00100000)
value POINTER_FLAG_INCONTACT (0x00000004)
value POINTER_FLAG_INRANGE (0x00000002)
value POINTER_FLAG_NEW (0x00000001)
value POINTER_FLAG_NONE (0x00000000)
value POINTER_FLAG_PRIMARY (0x00002000)
value POINTER_FLAG_SECONDBUTTON (0x00000020)
value POINTER_FLAG_THIRDBUTTON (0x00000040)
value POINTER_FLAG_UP (0x00040000)
value POINTER_FLAG_UPDATE (0x00020000)
value POINTER_FLAG_WHEEL (0x00080000)
value POINTER_MESSAGE_FLAG_CANCELED (0x00008000)
value POINTER_MESSAGE_FLAG_CONFIDENCE (0x00004000)
value POINTER_MESSAGE_FLAG_FIFTHBUTTON (0x00000100)
value POINTER_MESSAGE_FLAG_FIRSTBUTTON (0x00000010)
value POINTER_MESSAGE_FLAG_FOURTHBUTTON (0x00000080)
value POINTER_MESSAGE_FLAG_INCONTACT (0x00000004)
value POINTER_MESSAGE_FLAG_INRANGE (0x00000002)
value POINTER_MESSAGE_FLAG_NEW (0x00000001)
value POINTER_MESSAGE_FLAG_PRIMARY (0x00002000)
value POINTER_MESSAGE_FLAG_SECONDBUTTON (0x00000020)
value POINTER_MESSAGE_FLAG_THIRDBUTTON (0x00000040)
value POINTER_MOD_CTRL ((0x0008))
value POINTER_MOD_SHIFT ((0x0004))
value POLICY_AUDIT_SUBCATEGORY_COUNT ((59))
value POLICY_SHOWREASONUI_ALWAYS (1)
value POLICY_SHOWREASONUI_NEVER (0)
value POLICY_SHOWREASONUI_SERVERONLY (3)
value POLICY_SHOWREASONUI_WORKSTATIONONLY (2)
value POLLERR (0x0001)
value POLLHUP (0x0002)
value POLLIN ((POLLRDNORM | POLLRDBAND))
value POLLNVAL (0x0004)
value POLLOUT ((POLLWRNORM))
value POLLPRI (0x0400)
value POLLRDBAND (0x0200)
value POLLRDNORM (0x0100)
value POLLWRBAND (0x0020)
value POLLWRNORM (0x0010)
value POLYFILL_LAST (2)
value POLYGONALCAPS (32)
value POPENCARDNAMEA_EX (POPENCARDNAME_EXA)
value POPENCARDNAMEW_EX (POPENCARDNAME_EXW)
value POPENCARDNAME_A (POPENCARDNAMEA)
value POPENCARDNAME_W (POPENCARDNAMEW)
value PORT_STATUS_DOOR_OPEN (7)
value PORT_STATUS_NO_TONER (6)
value PORT_STATUS_OFFLINE (1)
value PORT_STATUS_OUTPUT_BIN_FULL (4)
value PORT_STATUS_OUT_OF_MEMORY (9)
value PORT_STATUS_PAPER_JAM (2)
value PORT_STATUS_PAPER_OUT (3)
value PORT_STATUS_PAPER_PROBLEM (5)
value PORT_STATUS_POWER_SAVE (12)
value PORT_STATUS_TONER_LOW (10)
value PORT_STATUS_TYPE_ERROR (1)
value PORT_STATUS_TYPE_INFO (3)
value PORT_STATUS_TYPE_WARNING (2)
value PORT_STATUS_USER_INTERVENTION (8)
value PORT_STATUS_WARMING_UP (11)
value PORT_TYPE_NET_ATTACHED (0x0008)
value PORT_TYPE_READ (0x0002)
value PORT_TYPE_REDIRECTED (0x0004)
value PORT_TYPE_WRITE (0x0001)
value POSITIVE_INFINITY_RATE (0xFFFFFFFE)
value POSTSCRIPT_DATA (37)
value POSTSCRIPT_IDENTIFY (4117)
value POSTSCRIPT_IGNORE (38)
value POSTSCRIPT_INJECTION (4118)
value POSTSCRIPT_PASSTHROUGH (4115)
value POWERBUTTON_ACTION_INDEX_HIBERNATE (2)
value POWERBUTTON_ACTION_INDEX_NOTHING (0)
value POWERBUTTON_ACTION_INDEX_SHUTDOWN (3)
value POWERBUTTON_ACTION_INDEX_SLEEP (1)
value POWERBUTTON_ACTION_INDEX_TURN_OFF_THE_DISPLAY (4)
value POWERBUTTON_ACTION_VALUE_HIBERNATE (3)
value POWERBUTTON_ACTION_VALUE_NOTHING (0)
value POWERBUTTON_ACTION_VALUE_SHUTDOWN (6)
value POWERBUTTON_ACTION_VALUE_SLEEP (2)
value POWERBUTTON_ACTION_VALUE_TURN_OFF_THE_DISPLAY (8)
value POWER_ACTION_ACPI_CRITICAL (0x01000000)
value POWER_ACTION_ACPI_USER_NOTIFY (0x02000000)
value POWER_ACTION_CRITICAL (0x80000000)
value POWER_ACTION_DIRECTED_DRIPS (0x04000000)
value POWER_ACTION_DISABLE_WAKES (0x40000000)
value POWER_ACTION_DOZE_TO_HIBERNATE (0x00000020)
value POWER_ACTION_HIBERBOOT (0x00000008)
value POWER_ACTION_LIGHTEST_FIRST (0x10000000)
value POWER_ACTION_LOCK_CONSOLE (0x20000000)
value POWER_ACTION_OVERRIDE_APPS (0x00000004)
value POWER_ACTION_PSEUDO_TRANSITION (0x08000000)
value POWER_ACTION_QUERY_ALLOWED (0x00000001)
value POWER_ACTION_UI_ALLOWED (0x00000002)
value POWER_ACTION_USER_NOTIFY (0x00000010)
value POWER_CONNECTIVITY_IN_STANDBY_DISABLED (0)
value POWER_CONNECTIVITY_IN_STANDBY_ENABLED (1)
value POWER_CONNECTIVITY_IN_STANDBY_SYSTEM_MANAGED (2)
value POWER_DEVICE_IDLE_POLICY_CONSERVATIVE (1)
value POWER_DEVICE_IDLE_POLICY_PERFORMANCE (0)
value POWER_DISCONNECTED_STANDBY_MODE_AGGRESSIVE (1)
value POWER_DISCONNECTED_STANDBY_MODE_NORMAL (0)
value POWER_FORCE_TRIGGER_RESET (0x80000000)
value POWER_LEVEL_USER_NOTIFY_EXEC (0x00000004)
value POWER_LEVEL_USER_NOTIFY_SOUND (0x00000002)
value POWER_LEVEL_USER_NOTIFY_TEXT (0x00000001)
value POWER_PLATFORM_ROLE_VERSION (POWER_PLATFORM_ROLE_V2)
value POWER_PLATFORM_ROLE_VERSION_MAX (POWER_PLATFORM_ROLE_V2_MAX)
value POWER_REQUEST_CONTEXT_DETAILED_STRING (DIAGNOSTIC_REASON_DETAILED_STRING)
value POWER_REQUEST_CONTEXT_SIMPLE_STRING (DIAGNOSTIC_REASON_SIMPLE_STRING)
value POWER_REQUEST_CONTEXT_VERSION (DIAGNOSTIC_REASON_VERSION)
value POWER_SETTING_VALUE_VERSION ((0x1))
value POWER_SYSTEM_MAXIMUM (7)
value POWER_USER_NOTIFY_BUTTON (0x00000008)
value POWER_USER_NOTIFY_FORCED_SHUTDOWN (0x00000020)
value POWER_USER_NOTIFY_SHUTDOWN (0x00000010)
value PO_DELETE (0x0013)
value PO_PORTCHANGE (0x0020)
value PO_RENAME (0x0014)
value PO_REN_PORT (0x0034)
value PO_THROTTLE_ADAPTIVE (3)
value PO_THROTTLE_CONSTANT (1)
value PO_THROTTLE_DEGRADE (2)
value PO_THROTTLE_MAXIMUM (4)
value PO_THROTTLE_NONE (0)
value PPCAPS_BOOKLET_EDGE (( 0x00000001 ))
value PPCAPS_BORDER_PRINT (( 0x00000001 ))
value PPCAPS_REVERSE_PAGES_FOR_REVERSE_DUPLEX (( 0x00000001 ))
value PPCAPS_RIGHT_THEN_DOWN (( 0x00000001 ))
value PPCAPS_SQUARE_SCALING (( 0x00000001 ))
value PPM_FIRMWARE_CPC (0x00040000)
value PPM_FIRMWARE_CSD (0x00000010)
value PPM_FIRMWARE_CST (0x00000008)
value PPM_FIRMWARE_LPI (0x00080000)
value PPM_FIRMWARE_OSC (0x00010000)
value PPM_FIRMWARE_PCCH (0x00004000)
value PPM_FIRMWARE_PCCP (0x00008000)
value PPM_FIRMWARE_PCT (0x00000020)
value PPM_FIRMWARE_PDC (0x00020000)
value PPM_FIRMWARE_PPC (0x00000100)
value PPM_FIRMWARE_PSD (0x00000200)
value PPM_FIRMWARE_PSS (0x00000040)
value PPM_FIRMWARE_PTC (0x00000400)
value PPM_FIRMWARE_TPC (0x00001000)
value PPM_FIRMWARE_TSD (0x00002000)
value PPM_FIRMWARE_TSS (0x00000800)
value PPM_FIRMWARE_XPSS (0x00000080)
value PPM_IDLE_IMPLEMENTATION_CSTATES (0x00000001)
value PPM_IDLE_IMPLEMENTATION_LPISTATES (0x00000004)
value PPM_IDLE_IMPLEMENTATION_MICROPEP (0x00000003)
value PPM_IDLE_IMPLEMENTATION_NONE (0x00000000)
value PPM_IDLE_IMPLEMENTATION_PEP (0x00000002)
value PPM_PERFORMANCE_IMPLEMENTATION_CPPC (0x00000003)
value PPM_PERFORMANCE_IMPLEMENTATION_NONE (0x00000000)
value PPM_PERFORMANCE_IMPLEMENTATION_PEP (0x00000004)
value PPM_PERFORMANCE_IMPLEMENTATION_PSTATES (0x00000001)
value PP_ADMIN_PIN (31)
value PP_APPLI_CERT (18)
value PP_CERTCHAIN (9)
value PP_CHANGE_PASSWORD (7)
value PP_CLIENT_HWND (1)
value PP_CONTAINER (6)
value PP_CONTEXT_INFO (11)
value PP_CRYPT_COUNT_KEY_USE (41)
value PP_DELETEKEY (24)
value PP_DISMISS_PIN_UI_SEC (49)
value PP_ENUMALGS (1)
value PP_ENUMALGS_EX (22)
value PP_ENUMCONTAINERS (2)
value PP_ENUMELECTROOTS (26)
value PP_ENUMEX_SIGNING_PROT (40)
value PP_ENUMMANDROOTS (25)
value PP_IMPTYPE (3)
value PP_IS_PFX_EPHEMERAL (50)
value PP_KEYEXCHANGE_ALG (14)
value PP_KEYEXCHANGE_KEYSIZE (12)
value PP_KEYEXCHANGE_PIN (32)
value PP_KEYSET_SEC_DESCR (8)
value PP_KEYSET_TYPE (27)
value PP_KEYSPEC (39)
value PP_KEYSTORAGE (17)
value PP_KEYX_KEYSIZE_INC (35)
value PP_KEY_TYPE_SUBTYPE (10)
value PP_NAME (4)
value PP_PIN_PROMPT_STRING (44)
value PP_PROVTYPE (16)
value PP_ROOT_CERTSTORE (46)
value PP_SECURE_KEYEXCHANGE_PIN (47)
value PP_SECURE_SIGNATURE_PIN (48)
value PP_SESSION_KEYSIZE (20)
value PP_SGC_INFO (37)
value PP_SIGNATURE_ALG (15)
value PP_SIGNATURE_KEYSIZE (13)
value PP_SIGNATURE_PIN (33)
value PP_SIG_KEYSIZE_INC (34)
value PP_SMARTCARD_GUID (45)
value PP_SMARTCARD_READER (43)
value PP_SMARTCARD_READER_ICON (47)
value PP_SYM_KEYSIZE (19)
value PP_UI_PROMPT (21)
value PP_UNIQUE_CONTAINER (36)
value PP_USER_CERTSTORE (42)
value PP_USE_HARDWARE_RNG (38)
value PP_VERSION (5)
value PRAGMA_DEPRECATED_DDK (0)
value PRESENTATION_ERROR_LOST (_HRESULT_TYPEDEF_(0x88810001L))
value PRF_CHECKVISIBLE (0x00000001L)
value PRF_CHILDREN (0x00000010L)
value PRF_CLIENT (0x00000004L)
value PRF_ERASEBKGND (0x00000008L)
value PRF_NONCLIENT (0x00000002L)
value PRF_OWNED (0x00000020L)
value PRINTACTION_DOCUMENTDEFAULTS (6)
value PRINTACTION_NETINSTALL (2)
value PRINTACTION_NETINSTALLLINK (3)
value PRINTACTION_OPEN (0)
value PRINTACTION_OPENNETPRN (5)
value PRINTACTION_PROPERTIES (1)
value PRINTACTION_SERVERPROPERTIES (7)
value PRINTACTION_TESTPAGE (4)
value PRINTDLGEXORD (1549)
value PRINTDLGORD (1538)
value PRINTER_ACCESS_ADMINISTER (0x00000004)
value PRINTER_ACCESS_MANAGE_LIMITED (0x00000040)
value PRINTER_ACCESS_USE (0x00000008)
value PRINTER_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | PRINTER_ACCESS_ADMINISTER | PRINTER_ACCESS_USE))
value PRINTER_ATTRIBUTE_DEFAULT (0x00000004)
value PRINTER_ATTRIBUTE_DIRECT (0x00000002)
value PRINTER_ATTRIBUTE_DO_COMPLETE_FIRST (0x00000200)
value PRINTER_ATTRIBUTE_ENABLE_BIDI (0x00000800)
value PRINTER_ATTRIBUTE_ENABLE_DEVQ (0x00000080)
value PRINTER_ATTRIBUTE_ENTERPRISE_CLOUD (0x00800000)
value PRINTER_ATTRIBUTE_FAX (0x00004000)
value PRINTER_ATTRIBUTE_FRIENDLY_NAME (0x00100000)
value PRINTER_ATTRIBUTE_HIDDEN (0x00000020)
value PRINTER_ATTRIBUTE_KEEPPRINTEDJOBS (0x00000100)
value PRINTER_ATTRIBUTE_LOCAL (0x00000040)
value PRINTER_ATTRIBUTE_MACHINE (0x00080000)
value PRINTER_ATTRIBUTE_NETWORK (0x00000010)
value PRINTER_ATTRIBUTE_PER_USER (0x00400000)
value PRINTER_ATTRIBUTE_PUBLISHED (0x00002000)
value PRINTER_ATTRIBUTE_PUSHED_MACHINE (0x00040000)
value PRINTER_ATTRIBUTE_PUSHED_USER (0x00020000)
value PRINTER_ATTRIBUTE_QUEUED (0x00000001)
value PRINTER_ATTRIBUTE_RAW_ONLY (0x00001000)
value PRINTER_ATTRIBUTE_SHARED (0x00000008)
value PRINTER_ATTRIBUTE_TS (0x00008000)
value PRINTER_ATTRIBUTE_TS_GENERIC_DRIVER (0x00200000)
value PRINTER_ATTRIBUTE_WORK_OFFLINE (0x00000400)
value PRINTER_CHANGE_ADD_FORM (0x00010000)
value PRINTER_CHANGE_ADD_JOB (0x00000100)
value PRINTER_CHANGE_ADD_PORT (0x00100000)
value PRINTER_CHANGE_ADD_PRINTER (0x00000001)
value PRINTER_CHANGE_ADD_PRINTER_DRIVER (0x10000000)
value PRINTER_CHANGE_ADD_PRINT_PROCESSOR (0x01000000)
value PRINTER_CHANGE_ALL (0x7F77FFFF)
value PRINTER_CHANGE_CONFIGURE_PORT (0x00200000)
value PRINTER_CHANGE_DELETE_FORM (0x00040000)
value PRINTER_CHANGE_DELETE_JOB (0x00000400)
value PRINTER_CHANGE_DELETE_PORT (0x00400000)
value PRINTER_CHANGE_DELETE_PRINTER (0x00000004)
value PRINTER_CHANGE_DELETE_PRINTER_DRIVER (0x40000000)
value PRINTER_CHANGE_DELETE_PRINT_PROCESSOR (0x04000000)
value PRINTER_CHANGE_FAILED_CONNECTION_PRINTER (0x00000008)
value PRINTER_CHANGE_FORM (0x00070000)
value PRINTER_CHANGE_JOB (0x0000FF00)
value PRINTER_CHANGE_PORT (0x00700000)
value PRINTER_CHANGE_PRINTER (0x000000FF)
value PRINTER_CHANGE_PRINTER_DRIVER (0x70000000)
value PRINTER_CHANGE_PRINT_PROCESSOR (0x07000000)
value PRINTER_CHANGE_SERVER (0x08000000)
value PRINTER_CHANGE_SET_FORM (0x00020000)
value PRINTER_CHANGE_SET_JOB (0x00000200)
value PRINTER_CHANGE_SET_PRINTER (0x00000002)
value PRINTER_CHANGE_SET_PRINTER_DRIVER (0x20000000)
value PRINTER_CHANGE_TIMEOUT (0x80000000)
value PRINTER_CHANGE_WRITE_JOB (0x00000800)
value PRINTER_CONNECTION_MISMATCH (0x00000020)
value PRINTER_CONNECTION_NO_UI (0x00000040)
value PRINTER_CONTROL_PAUSE (1)
value PRINTER_CONTROL_PURGE (3)
value PRINTER_CONTROL_RESUME (2)
value PRINTER_CONTROL_SET_STATUS (4)
value PRINTER_DRIVER_CATEGORY_CLOUD (0x00002000)
value PRINTER_DRIVER_CATEGORY_FAX (0x00000040)
value PRINTER_DRIVER_CATEGORY_FILE (0x00000080)
value PRINTER_DRIVER_CATEGORY_SERVICE (0x00000200)
value PRINTER_DRIVER_CATEGORY_VIRTUAL (0x00000100)
value PRINTER_DRIVER_CLASS (0x00000008)
value PRINTER_DRIVER_DERIVED (0x00000010)
value PRINTER_DRIVER_NOT_SHAREABLE (0x00000020)
value PRINTER_DRIVER_PACKAGE_AWARE (0x00000001)
value PRINTER_DRIVER_SANDBOX_DISABLED (0x00000800)
value PRINTER_DRIVER_SANDBOX_ENABLED (0x00000004)
value PRINTER_DRIVER_SOFT_RESET_REQUIRED (0x00000400)
value PRINTER_DRIVER_XPS (0x00000002)
value PRINTER_ENUM_CATEGORY_ALL (0x02000000)
value PRINTER_ENUM_CONNECTIONS (0x00000004)
value PRINTER_ENUM_CONTAINER (0x00008000)
value PRINTER_ENUM_DEFAULT (0x00000001)
value PRINTER_ENUM_EXPAND (0x00004000)
value PRINTER_ENUM_FAVORITE (0x00000004)
value PRINTER_ENUM_HIDE (0x01000000)
value PRINTER_ENUM_ICONMASK (0x00ff0000)
value PRINTER_ENUM_LOCAL (0x00000002)
value PRINTER_ENUM_NAME (0x00000008)
value PRINTER_ENUM_NETWORK (0x00000040)
value PRINTER_ENUM_REMOTE (0x00000010)
value PRINTER_ENUM_SHARED (0x00000020)
value PRINTER_ERROR_INFORMATION (0x80000000)
value PRINTER_ERROR_JAM (0x00000002)
value PRINTER_ERROR_OUTOFPAPER (0x00000001)
value PRINTER_ERROR_OUTOFTONER (0x00000004)
value PRINTER_ERROR_SEVERE (0x20000000)
value PRINTER_ERROR_WARNING (0x40000000)
value PRINTER_EXECUTE ((STANDARD_RIGHTS_EXECUTE | PRINTER_ACCESS_USE))
value PRINTER_FONTTYPE (0x4000)
value PRINTER_NOTIFY_CATEGORY_ALL (0x001000)
value PRINTER_NOTIFY_FIELD_ATTRIBUTES (0x0D)
value PRINTER_NOTIFY_FIELD_AVERAGE_PPM (0x15)
value PRINTER_NOTIFY_FIELD_BRANCH_OFFICE_PRINTING (0x1C)
value PRINTER_NOTIFY_FIELD_BYTES_PRINTED (0x19)
value PRINTER_NOTIFY_FIELD_CJOBS (0x14)
value PRINTER_NOTIFY_FIELD_COMMENT (0x05)
value PRINTER_NOTIFY_FIELD_DATATYPE (0x0B)
value PRINTER_NOTIFY_FIELD_DEFAULT_PRIORITY (0x0F)
value PRINTER_NOTIFY_FIELD_DEVMODE (0x07)
value PRINTER_NOTIFY_FIELD_DRIVER_NAME (0x04)
value PRINTER_NOTIFY_FIELD_FRIENDLY_NAME (0x1B)
value PRINTER_NOTIFY_FIELD_LOCATION (0x06)
value PRINTER_NOTIFY_FIELD_OBJECT_GUID (0x1A)
value PRINTER_NOTIFY_FIELD_PAGES_PRINTED (0x17)
value PRINTER_NOTIFY_FIELD_PARAMETERS (0x0A)
value PRINTER_NOTIFY_FIELD_PORT_NAME (0x03)
value PRINTER_NOTIFY_FIELD_PRINTER_NAME (0x01)
value PRINTER_NOTIFY_FIELD_PRINT_PROCESSOR (0x09)
value PRINTER_NOTIFY_FIELD_PRIORITY (0x0E)
value PRINTER_NOTIFY_FIELD_SECURITY_DESCRIPTOR (0x0C)
value PRINTER_NOTIFY_FIELD_SEPFILE (0x08)
value PRINTER_NOTIFY_FIELD_SERVER_NAME (0x00)
value PRINTER_NOTIFY_FIELD_SHARE_NAME (0x02)
value PRINTER_NOTIFY_FIELD_START_TIME (0x10)
value PRINTER_NOTIFY_FIELD_STATUS (0x12)
value PRINTER_NOTIFY_FIELD_STATUS_STRING (0x13)
value PRINTER_NOTIFY_FIELD_TOTAL_BYTES (0x18)
value PRINTER_NOTIFY_FIELD_TOTAL_PAGES (0x16)
value PRINTER_NOTIFY_FIELD_UNTIL_TIME (0x11)
value PRINTER_NOTIFY_INFO_DISCARDED (0x01)
value PRINTER_NOTIFY_OPTIONS_REFRESH (0x01)
value PRINTER_NOTIFY_TYPE (0x00)
value PRINTER_READ ((STANDARD_RIGHTS_READ | PRINTER_ACCESS_USE))
value PRINTER_STATUS_BUSY (0x00000200)
value PRINTER_STATUS_DOOR_OPEN (0x00400000)
value PRINTER_STATUS_DRIVER_UPDATE_NEEDED (0x04000000)
value PRINTER_STATUS_ERROR (0x00000002)
value PRINTER_STATUS_INITIALIZING (0x00008000)
value PRINTER_STATUS_IO_ACTIVE (0x00000100)
value PRINTER_STATUS_MANUAL_FEED (0x00000020)
value PRINTER_STATUS_NOT_AVAILABLE (0x00001000)
value PRINTER_STATUS_NO_TONER (0x00040000)
value PRINTER_STATUS_OFFLINE (0x00000080)
value PRINTER_STATUS_OUTPUT_BIN_FULL (0x00000800)
value PRINTER_STATUS_OUT_OF_MEMORY (0x00200000)
value PRINTER_STATUS_PAGE_PUNT (0x00080000)
value PRINTER_STATUS_PAPER_JAM (0x00000008)
value PRINTER_STATUS_PAPER_OUT (0x00000010)
value PRINTER_STATUS_PAPER_PROBLEM (0x00000040)
value PRINTER_STATUS_PAUSED (0x00000001)
value PRINTER_STATUS_PENDING_DELETION (0x00000004)
value PRINTER_STATUS_POWER_SAVE (0x01000000)
value PRINTER_STATUS_PRINTING (0x00000400)
value PRINTER_STATUS_PROCESSING (0x00004000)
value PRINTER_STATUS_SERVER_OFFLINE (0x02000000)
value PRINTER_STATUS_SERVER_UNKNOWN (0x00800000)
value PRINTER_STATUS_TONER_LOW (0x00020000)
value PRINTER_STATUS_USER_INTERVENTION (0x00100000)
value PRINTER_STATUS_WAITING (0x00002000)
value PRINTER_STATUS_WARMING_UP (0x00010000)
value PRINTER_WRITE ((STANDARD_RIGHTS_WRITE | PRINTER_ACCESS_USE))
value PRINTRATEUNIT_CPS (2)
value PRINTRATEUNIT_IPM (4)
value PRINTRATEUNIT_LPM (3)
value PRINTRATEUNIT_PPM (1)
value PRINT_PROP_FORCE_NAME (0x01)
value PRIVATEKEYBLOB (0x7)
value PRIVATE_NAMESPACE_FLAG_DESTROY (0x00000001)
value PRIVILEGE_SET_ALL_NECESSARY ((1))
value PRNSETUPDLGORD (1539)
value PROCESSOR_ARCHITECTURE_ALPHA (2)
value PROCESSOR_ARCHITECTURE_ARM (5)
value PROCESSOR_ARCHITECTURE_INTEL (0)
value PROCESSOR_ARCHITECTURE_MIPS (1)
value PROCESSOR_ARCHITECTURE_MSIL (8)
value PROCESSOR_ARCHITECTURE_NEUTRAL (11)
value PROCESSOR_ARCHITECTURE_PPC (3)
value PROCESSOR_ARCHITECTURE_SHX (4)
value PROCESSOR_ARCHITECTURE_UNKNOWN (0xFFFF)
value PROCESSOR_DUTY_CYCLING_DISABLED (0)
value PROCESSOR_DUTY_CYCLING_ENABLED (1)
value PROCESSOR_IDLESTATE_POLICY_COUNT (0x3)
value PROCESSOR_INTEL_PENTIUM (586)
value PROCESSOR_OPTIL (0x494f)
value PROCESSOR_PERF_AUTONOMOUS_MODE_DISABLED (0)
value PROCESSOR_PERF_AUTONOMOUS_MODE_ENABLED (1)
value PROCESSOR_PERF_BOOST_MODE_AGGRESSIVE (2)
value PROCESSOR_PERF_BOOST_MODE_AGGRESSIVE_AT_GUARANTEED (5)
value PROCESSOR_PERF_BOOST_MODE_DISABLED (0)
value PROCESSOR_PERF_BOOST_MODE_EFFICIENT_AGGRESSIVE (4)
value PROCESSOR_PERF_BOOST_MODE_EFFICIENT_AGGRESSIVE_AT_GUARANTEED (6)
value PROCESSOR_PERF_BOOST_MODE_EFFICIENT_ENABLED (3)
value PROCESSOR_PERF_BOOST_MODE_ENABLED (1)
value PROCESSOR_PERF_BOOST_MODE_MAX (PROCESSOR_PERF_BOOST_MODE_EFFICIENT_AGGRESSIVE_AT_GUARANTEED)
value PROCESSOR_PERF_BOOST_POLICY_DISABLED (0)
value PROCESSOR_PERF_BOOST_POLICY_MAX (100)
value PROCESSOR_PERF_ENERGY_PREFERENCE (0)
value PROCESSOR_PERF_MAXIMUM_ACTIVITY_WINDOW (1270000000)
value PROCESSOR_PERF_MINIMUM_ACTIVITY_WINDOW (0)
value PROCESSOR_PERF_PERFORMANCE_PREFERENCE (0xff)
value PROCESSOR_STRONGARM (2577)
value PROCESSOR_THROTTLE_AUTOMATIC (2)
value PROCESSOR_THROTTLE_DISABLED (0)
value PROCESSOR_THROTTLE_ENABLED (1)
value PROCESS_AFFINITY_ENABLE_AUTO_UPDATE (0x00000001UL)
value PROCESS_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | SYNCHRONIZE | 0xFFFF))
value PROCESS_CREATE_PROCESS ((0x0080))
value PROCESS_CREATE_THREAD ((0x0002))
value PROCESS_CREATION_ALL_APPLICATION_PACKAGES_OPT_OUT (0x01)
value PROCESS_CREATION_CHILD_PROCESS_OVERRIDE (0x02)
value PROCESS_CREATION_CHILD_PROCESS_RESTRICTED (0x01)
value PROCESS_CREATION_CHILD_PROCESS_RESTRICTED_UNLESS_SECURE (0x04)
value PROCESS_CREATION_DESKTOP_APP_BREAKAWAY_DISABLE_PROCESS_TREE (0x02)
value PROCESS_CREATION_DESKTOP_APP_BREAKAWAY_ENABLE_PROCESS_TREE (0x01)
value PROCESS_CREATION_DESKTOP_APP_BREAKAWAY_OVERRIDE (0x04)
value PROCESS_CREATION_MITIGATION_POLICY_DEP_ATL_THUNK_ENABLE (0x02)
value PROCESS_CREATION_MITIGATION_POLICY_DEP_ENABLE (0x01)
value PROCESS_CREATION_MITIGATION_POLICY_SEHOP_ENABLE (0x04)
value PROCESS_DEP_DISABLE_ATL_THUNK_EMULATION (0x00000002)
value PROCESS_DEP_ENABLE (0x00000001)
value PROCESS_DUP_HANDLE ((0x0040))
value PROCESS_HEAP_ENTRY_BUSY (0x0004)
value PROCESS_HEAP_ENTRY_DDESHARE (0x0020)
value PROCESS_HEAP_ENTRY_MOVEABLE (0x0010)
value PROCESS_HEAP_REGION (0x0001)
value PROCESS_HEAP_SEG_ALLOC (0x0008)
value PROCESS_HEAP_UNCOMMITTED_RANGE (0x0002)
value PROCESS_LEAP_SECOND_INFO_FLAG_ENABLE_SIXTY_SECOND (0x1)
value PROCESS_LEAP_SECOND_INFO_VALID_FLAGS ((PROCESS_LEAP_SECOND_INFO_FLAG_ENABLE_SIXTY_SECOND))
value PROCESS_MODE_BACKGROUND_BEGIN (0x00100000)
value PROCESS_MODE_BACKGROUND_END (0x00200000)
value PROCESS_NAME_NATIVE (0x00000001)
value PROCESS_POWER_THROTTLING_CURRENT_VERSION (1)
value PROCESS_POWER_THROTTLING_EXECUTION_SPEED (0x1)
value PROCESS_POWER_THROTTLING_IGNORE_TIMER_RESOLUTION (0x4)
value PROCESS_POWER_THROTTLING_VALID_FLAGS (((PROCESS_POWER_THROTTLING_EXECUTION_SPEED | PROCESS_POWER_THROTTLING_IGNORE_TIMER_RESOLUTION)))
value PROCESS_QUERY_INFORMATION ((0x0400))
value PROCESS_QUERY_LIMITED_INFORMATION ((0x1000))
value PROCESS_SET_INFORMATION ((0x0200))
value PROCESS_SET_LIMITED_INFORMATION ((0x2000))
value PROCESS_SET_QUOTA ((0x0100))
value PROCESS_SET_SESSIONID ((0x0004))
value PROCESS_SUSPEND_RESUME ((0x0800))
value PROCESS_TERMINATE ((0x0001))
value PROCESS_TRUST_LABEL_SECURITY_INFORMATION ((0x00000080L))
value PROCESS_VM_OPERATION ((0x0008))
value PROCESS_VM_READ ((0x0010))
value PROCESS_VM_WRITE ((0x0020))
value PROC_IDLE_BUCKET_COUNT (6)
value PROC_IDLE_BUCKET_COUNT_EX (16)
value PROC_THREAD_ATTRIBUTE_ADDITIVE (0x00040000)
value PROC_THREAD_ATTRIBUTE_INPUT (0x00020000)
value PROC_THREAD_ATTRIBUTE_NUMBER (0x0000FFFF)
value PROC_THREAD_ATTRIBUTE_REPLACE_VALUE (0x00000001)
value PROC_THREAD_ATTRIBUTE_THREAD (0x00010000)
value PRODUCT_AZURESTACKHCI_SERVER_CORE (0x00000196)
value PRODUCT_AZURE_NANO_SERVER (0x000000A9)
value PRODUCT_AZURE_SERVER_CLOUDHOST (0x000000C7)
value PRODUCT_AZURE_SERVER_CLOUDMOS (0x000000C8)
value PRODUCT_AZURE_SERVER_CORE (0x000000A8)
value PRODUCT_BUSINESS (0x00000006)
value PRODUCT_BUSINESS_N (0x00000010)
value PRODUCT_CLOUD (0x000000B2)
value PRODUCT_CLOUDE (0x000000B7)
value PRODUCT_CLOUDEDITION (0x000000CB)
value PRODUCT_CLOUDEDITIONN (0x000000CA)
value PRODUCT_CLOUDEN (0x000000BA)
value PRODUCT_CLOUDN (0x000000B3)
value PRODUCT_CLOUD_HOST_INFRASTRUCTURE_SERVER (0x0000007C)
value PRODUCT_CLOUD_STORAGE_SERVER (0x0000006E)
value PRODUCT_CLUSTER_SERVER (0x00000012)
value PRODUCT_CLUSTER_SERVER_V (0x00000040)
value PRODUCT_CONNECTED_CAR (0x00000075)
value PRODUCT_CORE (0x00000065)
value PRODUCT_CORE_ARM (0x00000061)
value PRODUCT_CORE_CONNECTED (0x0000006F)
value PRODUCT_CORE_CONNECTED_COUNTRYSPECIFIC (0x00000074)
value PRODUCT_CORE_CONNECTED_N (0x00000071)
value PRODUCT_CORE_CONNECTED_SINGLELANGUAGE (0x00000073)
value PRODUCT_CORE_COUNTRYSPECIFIC (0x00000063)
value PRODUCT_CORE_N (0x00000062)
value PRODUCT_CORE_SINGLELANGUAGE (0x00000064)
value PRODUCT_DATACENTER_A_SERVER_CORE (0x00000091)
value PRODUCT_DATACENTER_EVALUATION_SERVER (0x00000050)
value PRODUCT_DATACENTER_EVALUATION_SERVER_CORE (0x0000009F)
value PRODUCT_DATACENTER_NANO_SERVER (0x0000008F)
value PRODUCT_DATACENTER_SERVER (0x00000008)
value PRODUCT_DATACENTER_SERVER_AZURE_EDITION (0x00000197)
value PRODUCT_DATACENTER_SERVER_CORE (0x0000000C)
value PRODUCT_DATACENTER_SERVER_CORE_AZURE_EDITION (0x00000198)
value PRODUCT_DATACENTER_SERVER_CORE_V (0x00000027)
value PRODUCT_DATACENTER_SERVER_V (0x00000025)
value PRODUCT_DATACENTER_WS_SERVER_CORE (0x00000093)
value PRODUCT_EDUCATION (0x00000079)
value PRODUCT_EDUCATION_N (0x0000007A)
value PRODUCT_EMBEDDED (0x00000041)
value PRODUCT_EMBEDDED_A (0x00000058)
value PRODUCT_EMBEDDED_AUTOMOTIVE (0x00000055)
value PRODUCT_EMBEDDED_E (0x0000005A)
value PRODUCT_EMBEDDED_EVAL (0x0000006B)
value PRODUCT_EMBEDDED_E_EVAL (0x0000006C)
value PRODUCT_EMBEDDED_INDUSTRY (0x00000059)
value PRODUCT_EMBEDDED_INDUSTRY_A (0x00000056)
value PRODUCT_EMBEDDED_INDUSTRY_A_E (0x0000005C)
value PRODUCT_EMBEDDED_INDUSTRY_E (0x0000005B)
value PRODUCT_EMBEDDED_INDUSTRY_EVAL (0x00000069)
value PRODUCT_EMBEDDED_INDUSTRY_E_EVAL (0x0000006A)
value PRODUCT_ENTERPRISE (0x00000004)
value PRODUCT_ENTERPRISEG (0x000000AB)
value PRODUCT_ENTERPRISEGN (0x000000AC)
value PRODUCT_ENTERPRISE_E (0x00000046)
value PRODUCT_ENTERPRISE_EVALUATION (0x00000048)
value PRODUCT_ENTERPRISE_N (0x0000001B)
value PRODUCT_ENTERPRISE_N_EVALUATION (0x00000054)
value PRODUCT_ENTERPRISE_S (0x0000007D)
value PRODUCT_ENTERPRISE_SERVER (0x0000000A)
value PRODUCT_ENTERPRISE_SERVER_CORE (0x0000000E)
value PRODUCT_ENTERPRISE_SERVER_CORE_V (0x00000029)
value PRODUCT_ENTERPRISE_SERVER_V (0x00000026)
value PRODUCT_ENTERPRISE_SUBSCRIPTION (0x0000008C)
value PRODUCT_ENTERPRISE_SUBSCRIPTION_N (0x0000008D)
value PRODUCT_ENTERPRISE_S_EVALUATION (0x00000081)
value PRODUCT_ENTERPRISE_S_N (0x0000007E)
value PRODUCT_ENTERPRISE_S_N_EVALUATION (0x00000082)
value PRODUCT_ESSENTIALBUSINESS_SERVER_ADDL (0x0000003C)
value PRODUCT_ESSENTIALBUSINESS_SERVER_ADDLSVC (0x0000003E)
value PRODUCT_ESSENTIALBUSINESS_SERVER_MGMT (0x0000003B)
value PRODUCT_ESSENTIALBUSINESS_SERVER_MGMTSVC (0x0000003D)
value PRODUCT_HOLOGRAPHIC (0x00000087)
value PRODUCT_HOLOGRAPHIC_BUSINESS (0x00000088)
value PRODUCT_HOME_BASIC (0x00000002)
value PRODUCT_HOME_BASIC_E (0x00000043)
value PRODUCT_HOME_BASIC_N (0x00000005)
value PRODUCT_HOME_PREMIUM (0x00000003)
value PRODUCT_HOME_PREMIUM_E (0x00000044)
value PRODUCT_HOME_PREMIUM_N (0x0000001A)
value PRODUCT_HOME_PREMIUM_SERVER (0x00000022)
value PRODUCT_HOME_SERVER (0x00000013)
value PRODUCT_HUBOS (0x000000B4)
value PRODUCT_HYPERV (0x0000002A)
value PRODUCT_ID_LENGTH (16)
value PRODUCT_INDUSTRY_HANDHELD (0x00000076)
value PRODUCT_IOTEDGEOS (0x000000BB)
value PRODUCT_IOTENTERPRISE (0x000000BC)
value PRODUCT_IOTENTERPRISES (0x000000BF)
value PRODUCT_IOTOS (0x000000B9)
value PRODUCT_IOTUAP (0x0000007B)
value PRODUCT_LITE (0x000000BD)
value PRODUCT_MEDIUMBUSINESS_SERVER_MANAGEMENT (0x0000001E)
value PRODUCT_MEDIUMBUSINESS_SERVER_MESSAGING (0x00000020)
value PRODUCT_MEDIUMBUSINESS_SERVER_SECURITY (0x0000001F)
value PRODUCT_MULTIPOINT_PREMIUM_SERVER (0x0000004D)
value PRODUCT_MULTIPOINT_STANDARD_SERVER (0x0000004C)
value PRODUCT_NANO_SERVER (0x0000006D)
value PRODUCT_ONECOREUPDATEOS (0x000000B6)
value PRODUCT_PPI_PRO (0x00000077)
value PRODUCT_PROFESSIONAL (0x00000030)
value PRODUCT_PROFESSIONAL_E (0x00000045)
value PRODUCT_PROFESSIONAL_EMBEDDED (0x0000003A)
value PRODUCT_PROFESSIONAL_N (0x00000031)
value PRODUCT_PROFESSIONAL_S (0x0000007F)
value PRODUCT_PROFESSIONAL_STUDENT (0x00000070)
value PRODUCT_PROFESSIONAL_STUDENT_N (0x00000072)
value PRODUCT_PROFESSIONAL_S_N (0x00000080)
value PRODUCT_PROFESSIONAL_WMC (0x00000067)
value PRODUCT_PRO_CHINA (0x0000008B)
value PRODUCT_PRO_FOR_EDUCATION (0x000000A4)
value PRODUCT_PRO_FOR_EDUCATION_N (0x000000A5)
value PRODUCT_PRO_SINGLE_LANGUAGE (0x0000008A)
value PRODUCT_PRO_WORKSTATION (0x000000A1)
value PRODUCT_PRO_WORKSTATION_N (0x000000A2)
value PRODUCT_SB_SOLUTION_SERVER (0x00000032)
value PRODUCT_SB_SOLUTION_SERVER_EM (0x00000036)
value PRODUCT_SERVERRDSH (0x000000AF)
value PRODUCT_SERVER_FOR_SB_SOLUTIONS (0x00000033)
value PRODUCT_SERVER_FOR_SB_SOLUTIONS_EM (0x00000037)
value PRODUCT_SERVER_FOR_SMALLBUSINESS (0x00000018)
value PRODUCT_SERVER_FOR_SMALLBUSINESS_V (0x00000023)
value PRODUCT_SERVER_FOUNDATION (0x00000021)
value PRODUCT_SMALLBUSINESS_SERVER (0x00000009)
value PRODUCT_SMALLBUSINESS_SERVER_PREMIUM (0x00000019)
value PRODUCT_SMALLBUSINESS_SERVER_PREMIUM_CORE (0x0000003F)
value PRODUCT_SOLUTION_EMBEDDEDSERVER (0x00000038)
value PRODUCT_SOLUTION_EMBEDDEDSERVER_CORE (0x00000039)
value PRODUCT_STANDARD_A_SERVER_CORE (0x00000092)
value PRODUCT_STANDARD_EVALUATION_SERVER (0x0000004F)
value PRODUCT_STANDARD_EVALUATION_SERVER_CORE (0x000000A0)
value PRODUCT_STANDARD_NANO_SERVER (0x00000090)
value PRODUCT_STANDARD_SERVER (0x00000007)
value PRODUCT_STANDARD_SERVER_CORE (0x0000000D)
value PRODUCT_STANDARD_SERVER_CORE_V (0x00000028)
value PRODUCT_STANDARD_SERVER_SOLUTIONS (0x00000034)
value PRODUCT_STANDARD_SERVER_SOLUTIONS_CORE (0x00000035)
value PRODUCT_STANDARD_SERVER_V (0x00000024)
value PRODUCT_STANDARD_WS_SERVER_CORE (0x00000094)
value PRODUCT_STARTER (0x0000000B)
value PRODUCT_STARTER_E (0x00000042)
value PRODUCT_STARTER_N (0x0000002F)
value PRODUCT_STORAGE_ENTERPRISE_SERVER (0x00000017)
value PRODUCT_STORAGE_ENTERPRISE_SERVER_CORE (0x0000002E)
value PRODUCT_STORAGE_EXPRESS_SERVER (0x00000014)
value PRODUCT_STORAGE_EXPRESS_SERVER_CORE (0x0000002B)
value PRODUCT_STORAGE_STANDARD_EVALUATION_SERVER (0x00000060)
value PRODUCT_STORAGE_STANDARD_SERVER (0x00000015)
value PRODUCT_STORAGE_STANDARD_SERVER_CORE (0x0000002C)
value PRODUCT_STORAGE_WORKGROUP_EVALUATION_SERVER (0x0000005F)
value PRODUCT_STORAGE_WORKGROUP_SERVER (0x00000016)
value PRODUCT_STORAGE_WORKGROUP_SERVER_CORE (0x0000002D)
value PRODUCT_THINPC (0x00000057)
value PRODUCT_ULTIMATE (0x00000001)
value PRODUCT_ULTIMATE_E (0x00000047)
value PRODUCT_ULTIMATE_N (0x0000001C)
value PRODUCT_UNDEFINED (0x00000000)
value PRODUCT_UNLICENSED (0xABCDABCD)
value PRODUCT_UTILITY_VM (0x00000095)
value PRODUCT_WEB_SERVER (0x00000011)
value PRODUCT_WEB_SERVER_CORE (0x0000001D)
value PRODUCT_XBOX_DURANGOHOSTOS (0x000000C4)
value PRODUCT_XBOX_ERAOS (0x000000C3)
value PRODUCT_XBOX_GAMEOS (0x000000C2)
value PRODUCT_XBOX_KEYSTONE (0x000000C6)
value PRODUCT_XBOX_SCARLETTHOSTOS (0x000000C5)
value PRODUCT_XBOX_SYSTEMOS (0x000000C0)
value PROFILE_KERNEL (0x20000000)
value PROFILE_SERVER (0x40000000)
value PROFILE_USER (0x10000000)
value PROGRESS_CANCEL (1)
value PROGRESS_CONTINUE (0)
value PROGRESS_QUIET (3)
value PROGRESS_STOP (2)
value PROJFS_PROTOCOL_VERSION (3)
value PROOF_QUALITY (2)
value PROPSETFLAG_ANSI (( 2 ))
value PROPSETFLAG_CASE_SENSITIVE (( 8 ))
value PROPSETFLAG_DEFAULT (( 0 ))
value PROPSETFLAG_NONSIMPLE (( 1 ))
value PROPSETFLAG_UNBUFFERED (( 4 ))
value PROPSETHDR_OSVERSION_UNKNOWN (0xFFFFFFFF)
value PROPSET_BEHAVIOR_CASE_SENSITIVE (( 1 ))
value PROPSHEETHEADER (PROPSHEETHEADERA)
value PROPSHEETPAGE (PROPSHEETPAGEA)
value PROPSHEETPAGE_LATEST (PROPSHEETPAGEA_LATEST)
value PROP_LG_CXDLG (252)
value PROP_LG_CYDLG (218)
value PROP_MED_CXDLG (227)
value PROP_MED_CYDLG (215)
value PROP_SM_CXDLG (212)
value PROP_SM_CYDLG (188)
value PROTECTED_DACL_SECURITY_INFORMATION ((0x80000000L))
value PROTECTED_SACL_SECURITY_INFORMATION ((0x40000000L))
value PROTECTION_LEVEL_ANTIMALWARE_LIGHT (0x00000003)
value PROTECTION_LEVEL_AUTHENTICODE (0x00000007)
value PROTECTION_LEVEL_CODEGEN_LIGHT (0x00000006)
value PROTECTION_LEVEL_LSA_LIGHT (0x00000004)
value PROTECTION_LEVEL_NONE (0xFFFFFFFE)
value PROTECTION_LEVEL_PPL_APP (0x00000008)
value PROTECTION_LEVEL_SAME (0xFFFFFFFF)
value PROTECTION_LEVEL_WINDOWS (0x00000001)
value PROTECTION_LEVEL_WINDOWS_LIGHT (0x00000002)
value PROTECTION_LEVEL_WINTCB (0x00000005)
value PROTECTION_LEVEL_WINTCB_LIGHT (0x00000000)
value PROTOCOLFLAG_NO_PICS_CHECK (0x00000001)
value PROVIDER_KEEPS_VALUE_LENGTH (0x1)
value PROV_DH_SCHANNEL (18)
value PROV_DSS (3)
value PROV_DSS_DH (13)
value PROV_EC_ECDSA_FULL (16)
value PROV_EC_ECDSA_SIG (14)
value PROV_EC_ECNRA_FULL (17)
value PROV_EC_ECNRA_SIG (15)
value PROV_FORTEZZA (4)
value PROV_INTEL_SEC (22)
value PROV_MS_EXCHANGE (5)
value PROV_REPLACE_OWF (23)
value PROV_RNG (21)
value PROV_RSA_AES (24)
value PROV_RSA_FULL (1)
value PROV_RSA_SCHANNEL (12)
value PROV_RSA_SIG (2)
value PROV_SPYRUS_LYNKS (20)
value PROV_SSL (6)
value PRPC_ENDPOINT_TEMPLATE (PRPC_ENDPOINT_TEMPLATEA)
value PRPC_HTTP_TRANSPORT_CREDENTIALS (PRPC_HTTP_TRANSPORT_CREDENTIALS_A)
value PRPC_INTERFACE_TEMPLATE (PRPC_INTERFACE_TEMPLATEA)
value PRSPEC_LPWSTR (( 0 ))
value PRSPEC_PROPID (( 1 ))
value PR_JOBSTATUS (0x0000)
value PSBTN_APPLYNOW (4)
value PSBTN_BACK (0)
value PSBTN_CANCEL (5)
value PSBTN_FINISH (2)
value PSBTN_HELP (6)
value PSBTN_MAX (6)
value PSBTN_NEXT (1)
value PSBTN_OK (3)
value PSCARD_READERSTATE_A (PSCARD_READERSTATEA)
value PSCARD_READERSTATE_W (PSCARD_READERSTATEW)
value PSCB_BUTTONPRESSED (3)
value PSCB_INITIALIZED (1)
value PSCB_PRECREATE (2)
value PSD_DEFAULTMINMARGINS (0x00000000)
value PSD_DISABLEMARGINS (0x00000010)
value PSD_DISABLEORIENTATION (0x00000100)
value PSD_DISABLEPAGEPAINTING (0x00080000)
value PSD_DISABLEPAPER (0x00000200)
value PSD_DISABLEPRINTER (0x00000020)
value PSD_ENABLEPAGEPAINTHOOK (0x00040000)
value PSD_ENABLEPAGESETUPHOOK (0x00002000)
value PSD_ENABLEPAGESETUPTEMPLATE (0x00008000)
value PSD_ENABLEPAGESETUPTEMPLATEHANDLE (0x00020000)
value PSD_INHUNDREDTHSOFMILLIMETERS (0x00000008)
value PSD_INTHOUSANDTHSOFINCHES (0x00000004)
value PSD_INWININIINTLMEASURE (0x00000000)
value PSD_MARGINS (0x00000002)
value PSD_MINMARGINS (0x00000001)
value PSD_NONETWORKBUTTON (0x00200000)
value PSD_NOWARNING (0x00000080)
value PSD_RETURNDEFAULT (0x00000400)
value PSD_SHOWHELP (0x00000800)
value PSEC_WINNT_AUTH_IDENTITY (PSEC_WINNT_AUTH_IDENTITY_A)
value PSEUDOCONSOLE_INHERIT_CURSOR ((0x1))
value PSH_AEROWIZARD (0x00004000)
value PSH_DEFAULT (0x00000000)
value PSH_HASHELP (0x00000200)
value PSH_HEADER (0x00080000)
value PSH_HEADERBITMAP (0x08000000)
value PSH_MODELESS (0x00000400)
value PSH_NOAPPLYNOW (0x00000080)
value PSH_NOCONTEXTHELP (0x02000000)
value PSH_NOMARGIN (0x10000000)
value PSH_PROPSHEETPAGE (0x00000008)
value PSH_PROPTITLE (0x00000001)
value PSH_RESIZABLE (0x04000000)
value PSH_RTLREADING (0x00000800)
value PSH_STRETCHWATERMARK (0x00040000)
value PSH_USECALLBACK (0x00000100)
value PSH_USEHBMHEADER (0x00100000)
value PSH_USEHBMWATERMARK (0x00010000)
value PSH_USEHICON (0x00000002)
value PSH_USEHPLWATERMARK (0x00020000)
value PSH_USEICONID (0x00000004)
value PSH_USEPAGELANG (0x00200000)
value PSH_USEPSTARTPAGE (0x00000040)
value PSH_WATERMARK (0x00008000)
value PSH_WIZARD (0x00000020)
value PSH_WIZARDCONTEXTHELP (0x00001000)
value PSH_WIZARDHASFINISH (0x00000010)
value PSH_WIZARD_LITE (0x00400000)
value PSIDENT_GDICENTRIC (0)
value PSIDENT_PSCENTRIC (1)
value PSINJECT_BEGINDEFAULTS (12)
value PSINJECT_BEGINPAGESETUP (101)
value PSINJECT_BEGINPROLOG (14)
value PSINJECT_BEGINSETUP (16)
value PSINJECT_BEGINSTREAM (1)
value PSINJECT_BOUNDINGBOX (9)
value PSINJECT_COMMENTS (11)
value PSINJECT_DLFONT (0xdddddddd)
value PSINJECT_DOCNEEDEDRES (5)
value PSINJECT_DOCSUPPLIEDRES (6)
value PSINJECT_DOCUMENTPROCESSCOLORS (10)
value PSINJECT_DOCUMENTPROCESSCOLORSATEND (21)
value PSINJECT_ENDDEFAULTS (13)
value PSINJECT_ENDPAGECOMMENTS (107)
value PSINJECT_ENDPAGESETUP (102)
value PSINJECT_ENDPROLOG (15)
value PSINJECT_ENDSETUP (17)
value PSINJECT_ENDSTREAM (20)
value PSINJECT_EOF (19)
value PSINJECT_ORIENTATION (8)
value PSINJECT_PAGEBBOX (106)
value PSINJECT_PAGENUMBER (100)
value PSINJECT_PAGEORDER (7)
value PSINJECT_PAGES (4)
value PSINJECT_PAGESATEND (3)
value PSINJECT_PAGETRAILER (103)
value PSINJECT_PLATECOLOR (104)
value PSINJECT_PSADOBE (2)
value PSINJECT_SHOWPAGE (105)
value PSINJECT_TRAILER (18)
value PSINJECT_VMRESTORE (201)
value PSINJECT_VMSAVE (200)
value PSM_ADDPAGE ((WM_USER + 103))
value PSM_APPLY ((WM_USER + 110))
value PSM_CANCELTOCLOSE ((WM_USER + 107))
value PSM_CHANGED ((WM_USER + 104))
value PSM_ENABLEWIZBUTTONS ((WM_USER + 139))
value PSM_GETCURRENTPAGEHWND ((WM_USER + 118))
value PSM_GETRESULT ((WM_USER + 135))
value PSM_GETTABCONTROL ((WM_USER + 116))
value PSM_HWNDTOINDEX ((WM_USER + 129))
value PSM_IDTOINDEX ((WM_USER + 133))
value PSM_INDEXTOHWND ((WM_USER + 130))
value PSM_INDEXTOID ((WM_USER + 134))
value PSM_INDEXTOPAGE ((WM_USER + 132))
value PSM_INSERTPAGE ((WM_USER + 119))
value PSM_ISDIALOGMESSAGE ((WM_USER + 117))
value PSM_PAGETOINDEX ((WM_USER + 131))
value PSM_PRESSBUTTON ((WM_USER + 113))
value PSM_QUERYSIBLINGS ((WM_USER + 108))
value PSM_REBOOTSYSTEM ((WM_USER + 106))
value PSM_RECALCPAGESIZES ((WM_USER + 136))
value PSM_REMOVEPAGE ((WM_USER + 102))
value PSM_RESTARTWINDOWS ((WM_USER + 105))
value PSM_SETBUTTONTEXT (PSM_SETBUTTONTEXTW)
value PSM_SETBUTTONTEXTW ((WM_USER + 140))
value PSM_SETCURSEL ((WM_USER + 101))
value PSM_SETCURSELID ((WM_USER + 114))
value PSM_SETFINISHTEXT (PSM_SETFINISHTEXTA)
value PSM_SETFINISHTEXTA ((WM_USER + 115))
value PSM_SETFINISHTEXTW ((WM_USER + 121))
value PSM_SETHEADERSUBTITLE (PSM_SETHEADERSUBTITLEA)
value PSM_SETHEADERSUBTITLEA ((WM_USER + 127))
value PSM_SETHEADERSUBTITLEW ((WM_USER + 128))
value PSM_SETHEADERTITLE (PSM_SETHEADERTITLEA)
value PSM_SETHEADERTITLEA ((WM_USER + 125))
value PSM_SETHEADERTITLEW ((WM_USER + 126))
value PSM_SETNEXTTEXT (PSM_SETNEXTTEXTW)
value PSM_SETNEXTTEXTW ((WM_USER + 137))
value PSM_SETTITLE (PSM_SETTITLEA)
value PSM_SETTITLEA ((WM_USER + 111))
value PSM_SETTITLEW ((WM_USER + 120))
value PSM_SETWIZBUTTONS ((WM_USER + 112))
value PSM_SHOWWIZBUTTONS ((WM_USER + 138))
value PSM_UNCHANGED ((WM_USER + 109))
value PSNRET_INVALID (1)
value PSNRET_INVALID_NOCHANGEPAGE (2)
value PSNRET_MESSAGEHANDLED (3)
value PSNRET_NOERROR (0)
value PSN_APPLY ((PSN_FIRST-2))
value PSN_FIRST ((0U-200U))
value PSN_GETOBJECT ((PSN_FIRST-10))
value PSN_HELP ((PSN_FIRST-5))
value PSN_KILLACTIVE ((PSN_FIRST-1))
value PSN_LAST ((0U-299U))
value PSN_QUERYCANCEL ((PSN_FIRST-9))
value PSN_QUERYINITIALFOCUS ((PSN_FIRST-13))
value PSN_RESET ((PSN_FIRST-3))
value PSN_SETACTIVE ((PSN_FIRST-0))
value PSN_TRANSLATEACCELERATOR ((PSN_FIRST-12))
value PSN_WIZBACK ((PSN_FIRST-6))
value PSN_WIZFINISH ((PSN_FIRST-8))
value PSN_WIZNEXT ((PSN_FIRST-7))
value PSPCB_ADDREF (0)
value PSPCB_CREATE (2)
value PSPCB_RELEASE (1)
value PSPROTOCOL_ASCII (0)
value PSPROTOCOL_BCP (1)
value PSPROTOCOL_BINARY (3)
value PSPROTOCOL_TBCP (2)
value PSP_DEFAULT (0x00000000)
value PSP_DLGINDIRECT (0x00000001)
value PSP_HASHELP (0x00000020)
value PSP_HIDEHEADER (0x00000800)
value PSP_PREMATURE (0x00000400)
value PSP_RTLREADING (0x00000010)
value PSP_USECALLBACK (0x00000080)
value PSP_USEFUSIONCONTEXT (0x00004000)
value PSP_USEHEADERSUBTITLE (0x00002000)
value PSP_USEHEADERTITLE (0x00001000)
value PSP_USEHICON (0x00000002)
value PSP_USEICONID (0x00000004)
value PSP_USEREFPARENT (0x00000040)
value PSP_USETITLE (0x00000008)
value PST_FAX (((DWORD)0x00000021))
value PST_LAT (((DWORD)0x00000101))
value PST_MODEM (((DWORD)0x00000006))
value PST_NETWORK_BRIDGE (((DWORD)0x00000100))
value PST_PARALLELPORT (((DWORD)0x00000002))
value PST_SCANNER (((DWORD)0x00000022))
value PST_TCPIP_TELNET (((DWORD)0x00000102))
value PST_UNSPECIFIED (((DWORD)0x00000000))
value PSWIZBF_ELEVATIONREQUIRED (0x00000001)
value PSWIZB_BACK (0x00000001)
value PSWIZB_CANCEL (0x00000010)
value PSWIZB_DISABLEDFINISH (0x00000008)
value PSWIZB_FINISH (0x00000004)
value PSWIZB_NEXT (0x00000002)
value PSWIZB_RESTORE (1)
value PSWIZB_SHOW (0)
value PSWIZF_SETCOLOR (((UINT)(-1)))
value PS_ALTERNATE (8)
value PS_COSMETIC (0x00000000)
value PS_DASH (1)
value PS_DASHDOT (3)
value PS_DASHDOTDOT (4)
value PS_DOT (2)
value PS_ENDCAP_FLAT (0x00000200)
value PS_ENDCAP_MASK (0x00000F00)
value PS_ENDCAP_ROUND (0x00000000)
value PS_ENDCAP_SQUARE (0x00000100)
value PS_GEOMETRIC (0x00010000)
value PS_INSIDEFRAME (6)
value PS_JOIN_BEVEL (0x00001000)
value PS_JOIN_MASK (0x0000F000)
value PS_JOIN_MITER (0x00002000)
value PS_JOIN_ROUND (0x00000000)
value PS_NULL (5)
value PS_OPENTYPE_FONTTYPE (0x10000)
value PS_SOLID (0)
value PS_STYLE_MASK (0x0000000F)
value PS_TYPE_MASK (0x000F0000)
value PS_USERSTYLE (7)
value PT_BEZIERTO (0x04)
value PT_CLOSEFIGURE (0x01)
value PT_LINETO (0x02)
value PT_MOVETO (0x06)
value PUBLICKEYBLOB (0x6)
value PUBLICKEYBLOBEX (0xA)
value PURGE_RXABORT (0x0002)
value PURGE_RXCLEAR (0x0008)
value PURGE_TXABORT (0x0001)
value PURGE_TXCLEAR (0x0004)
value PVD_CONFIG (0x3001)
value PWR_CRITICALRESUME (3)
value PWR_FAIL ((-1))
value PWR_OK (1)
value PWR_SUSPENDREQUEST (1)
value PWR_SUSPENDRESUME (2)
value PW_CLIENTONLY (0x00000001)
value PW_RENDERFULLCONTENT (0x00000002)
value QDC_ALL_PATHS (0x00000001)
value QDC_DATABASE_CURRENT (0x00000004)
value QDC_INCLUDE_HMD (0x00000020)
value QDC_ONLY_ACTIVE_PATHS (0x00000002)
value QDC_VIRTUAL_MODE_AWARE (0x00000010)
value QDC_VIRTUAL_REFRESH_RATE_AWARE (0x00000040)
value QDI_DIBTOSCREEN (4)
value QDI_GETDIBITS (2)
value QDI_SETDIBITS (1)
value QDI_STRETCHDIB (8)
value QID_SYNC (0xFFFFFFFF)
value QOS_GENERAL_ID_BASE (2000)
value QOS_NOT_SPECIFIED (0xFFFFFFFF)
value QOS_OBJECT_DESTADDR ((0x00000004 + QOS_GENERAL_ID_BASE))
value QOS_OBJECT_END_OF_LIST ((0x00000001 + QOS_GENERAL_ID_BASE))
value QOS_OBJECT_SD_MODE ((0x00000002 + QOS_GENERAL_ID_BASE))
value QOS_OBJECT_SHAPING_RATE ((0x00000003 + QOS_GENERAL_ID_BASE))
value QS_ALLEVENTS ((QS_INPUT | QS_POSTMESSAGE | QS_TIMER | QS_PAINT | QS_HOTKEY))
value QS_ALLINPUT ((QS_INPUT | QS_POSTMESSAGE | QS_TIMER | QS_PAINT | QS_HOTKEY | QS_SENDMESSAGE))
value QS_ALLPOSTMESSAGE (0x0100)
value QS_HOTKEY (0x0080)
value QS_INPUT ((QS_MOUSE | QS_KEY | QS_RAWINPUT | QS_TOUCH | QS_POINTER))
value QS_KEY (0x0001)
value QS_MOUSE ((QS_MOUSEMOVE | QS_MOUSEBUTTON))
value QS_MOUSEBUTTON (0x0004)
value QS_MOUSEMOVE (0x0002)
value QS_PAINT (0x0020)
value QS_POINTER (0x1000)
value QS_POSTMESSAGE (0x0008)
value QS_RAWINPUT (0x0400)
value QS_SENDMESSAGE (0x0040)
value QS_TIMER (0x0010)
value QS_TOUCH (0x0800)
value QUERYDIBSUPPORT (3073)
value QUERYESCSUPPORT (8)
value QUERYROPSUPPORT (40)
value QUERY_ACTCTX_FLAG_ACTCTX_IS_ADDRESS ((0x00000010))
value QUERY_ACTCTX_FLAG_ACTCTX_IS_HMODULE ((0x00000008))
value QUERY_ACTCTX_FLAG_NO_ADDREF ((0x80000000))
value QUERY_ACTCTX_FLAG_USE_ACTIVE_ACTCTX ((0x00000004))
value QUERY_DEPENDENT_VOLUME_REQUEST_FLAG_GUEST_VOLUMES (0x2)
value QUERY_DEPENDENT_VOLUME_REQUEST_FLAG_HOST_VOLUMES (0x1)
value QUERY_FILE_LAYOUT_INCLUDE_EXTENTS ((0x00000008))
value QUERY_FILE_LAYOUT_INCLUDE_EXTRA_INFO ((0x00000010))
value QUERY_FILE_LAYOUT_INCLUDE_FILES_WITH_DSC_ATTRIBUTE ((0x00001000))
value QUERY_FILE_LAYOUT_INCLUDE_FULL_PATH_IN_NAMES ((0x00000040))
value QUERY_FILE_LAYOUT_INCLUDE_NAMES ((0x00000002))
value QUERY_FILE_LAYOUT_INCLUDE_ONLY_FILES_WITH_SPECIFIC_ATTRIBUTES ((0x00000800))
value QUERY_FILE_LAYOUT_INCLUDE_STREAMS ((0x00000004))
value QUERY_FILE_LAYOUT_INCLUDE_STREAMS_WITH_NO_CLUSTERS_ALLOCATED ((0x00000020))
value QUERY_FILE_LAYOUT_INCLUDE_STREAM_INFORMATION ((0x00000080))
value QUERY_FILE_LAYOUT_INCLUDE_STREAM_INFORMATION_FOR_DATA_ATTRIBUTE ((0x00002000))
value QUERY_FILE_LAYOUT_INCLUDE_STREAM_INFORMATION_FOR_DSC_ATTRIBUTE ((0x00000100))
value QUERY_FILE_LAYOUT_INCLUDE_STREAM_INFORMATION_FOR_EA_ATTRIBUTE ((0x00008000))
value QUERY_FILE_LAYOUT_INCLUDE_STREAM_INFORMATION_FOR_EFS_ATTRIBUTE ((0x00000400))
value QUERY_FILE_LAYOUT_INCLUDE_STREAM_INFORMATION_FOR_REPARSE_ATTRIBUTE ((0x00004000))
value QUERY_FILE_LAYOUT_INCLUDE_STREAM_INFORMATION_FOR_TXF_ATTRIBUTE ((0x00000200))
value QUERY_FILE_LAYOUT_REPARSE_DATA_INVALID ((0x0001))
value QUERY_FILE_LAYOUT_REPARSE_TAG_INVALID ((0x0002))
value QUERY_FILE_LAYOUT_RESTART ((0x00000001))
value QUERY_FILE_LAYOUT_SINGLE_INSTANCED ((0x00000001))
value QUERY_STORAGE_CLASSES_FLAGS_MEASURE_READ (0x40000000)
value QUERY_STORAGE_CLASSES_FLAGS_MEASURE_WRITE (0x80000000)
value QUERY_STORAGE_CLASSES_FLAGS_NO_DEFRAG_VOLUME (0x20000000)
value QUOTA_LIMITS_HARDWS_MAX_DISABLE (0x00000008)
value QUOTA_LIMITS_HARDWS_MAX_ENABLE (0x00000004)
value QUOTA_LIMITS_HARDWS_MIN_DISABLE (0x00000002)
value QUOTA_LIMITS_HARDWS_MIN_ENABLE (0x00000001)
value QUOTA_LIMITS_USE_DEFAULT_LIMITS (0x00000010)
value RANDOM_PADDING (2)
value RAND_MAX (0x7fff)
value RASTERCAPS (38)
value RASTER_FONTTYPE (0x0001)
value RC_BANDING (2)
value RC_BIGFONT (0x0400)
value RC_BITBLT (1)
value RC_DEVBITS (0x8000)
value RC_DIBTODEV (0x0200)
value RC_DI_BITMAP (0x0080)
value RC_FLOODFILL (0x1000)
value RC_OP_DX_OUTPUT (0x4000)
value RC_PALETTE (0x0100)
value RC_SAVEBITMAP (0x0040)
value RC_SCALING (4)
value RC_STRETCHBLT (0x0800)
value RC_STRETCHDIB (0x2000)
value RDH_RECTANGLES (1)
value RDW_ALLCHILDREN (0x0080)
value RDW_ERASE (0x0004)
value RDW_ERASENOW (0x0200)
value RDW_FRAME (0x0400)
value RDW_INTERNALPAINT (0x0002)
value RDW_INVALIDATE (0x0001)
value RDW_NOCHILDREN (0x0040)
value RDW_NOERASE (0x0020)
value RDW_NOFRAME (0x0800)
value RDW_NOINTERNALPAINT (0x0010)
value RDW_UPDATENOW (0x0100)
value RDW_VALIDATE (0x0008)
value READ_ATTRIBUTES (0xD0)
value READ_ATTRIBUTE_BUFFER_SIZE (512)
value READ_COMPRESSION_INFO_VALID (0x00000020)
value READ_CONTROL ((0x00020000L))
value READ_COPY_NUMBER_BYPASS_CACHE_FLAG (0x00000100)
value READ_COPY_NUMBER_KEY (0x52434e00)
value READ_THREAD_PROFILING_FLAG_DISPATCHING (0x00000001)
value READ_THREAD_PROFILING_FLAG_HARDWARE_COUNTERS (0x00000002)
value READ_THRESHOLDS (0xD1)
value READ_THRESHOLD_BUFFER_SIZE (512)
value REALTIME_PRIORITY_CLASS (0x00000100)
value REASON_HWINSTALL ((SHTDN_REASON_MAJOR_HARDWARE|SHTDN_REASON_MINOR_INSTALLATION))
value REASON_LEGACY_API (SHTDN_REASON_LEGACY_API)
value REASON_OTHER ((SHTDN_REASON_MAJOR_OTHER|SHTDN_REASON_MINOR_OTHER))
value REASON_PLANNED_FLAG (SHTDN_REASON_FLAG_PLANNED)
value REASON_SERVICEHANG ((SHTDN_REASON_MAJOR_SOFTWARE|SHTDN_REASON_MINOR_HUNG))
value REASON_SWHWRECONF ((SHTDN_REASON_MAJOR_SOFTWARE|SHTDN_REASON_MINOR_RECONFIG))
value REASON_SWINSTALL ((SHTDN_REASON_MAJOR_SOFTWARE|SHTDN_REASON_MINOR_INSTALLATION))
value REASON_UNKNOWN (SHTDN_REASON_UNKNOWN)
value REASON_UNSTABLE ((SHTDN_REASON_MAJOR_SYSTEM|SHTDN_REASON_MINOR_UNSTABLE))
value RECOVERED_READS_VALID (0x00000004)
value RECOVERED_WRITES_VALID (0x00000001)
value RECOVERY_DEFAULT_PING_INTERVAL (5000)
value REFERENCE_BLACK_MAX ((WORD)4000)
value REFERENCE_BLACK_MIN ((WORD)0)
value REFERENCE_WHITE_MAX ((WORD)10000)
value REFERENCE_WHITE_MIN ((WORD)6000)
value REGDB_E_BADTHREADINGMODEL (_HRESULT_TYPEDEF_(0x80040156L))
value REGDB_E_CLASSNOTREG (_HRESULT_TYPEDEF_(0x80040154L))
value REGDB_E_FIRST (0x80040150L)
value REGDB_E_IIDNOTREG (_HRESULT_TYPEDEF_(0x80040155L))
value REGDB_E_INVALIDVALUE (_HRESULT_TYPEDEF_(0x80040153L))
value REGDB_E_KEYMISSING (_HRESULT_TYPEDEF_(0x80040152L))
value REGDB_E_LAST (0x8004015FL)
value REGDB_E_PACKAGEPOLICYVIOLATION (_HRESULT_TYPEDEF_(0x80040157L))
value REGDB_E_READREGDB (_HRESULT_TYPEDEF_(0x80040150L))
value REGDB_E_WRITEREGDB (_HRESULT_TYPEDEF_(0x80040151L))
value REGDB_S_FIRST (0x00040150L)
value REGDB_S_LAST (0x0004015FL)
value REGISTERED (0x04)
value REGISTERING (0x00)
value REGISTERWORDENUMPROC (REGISTERWORDENUMPROCA)
value REGULAR_FONTTYPE (0x0400)
value REG_APP_HIVE ((0x00000010L))
value REG_APP_HIVE_OPEN_READ_ONLY ((REG_OPEN_READ_ONLY))
value REG_BOOT_HIVE ((0x00000400L))
value REG_CREATED_NEW_KEY ((0x00000001L))
value REG_FLUSH_HIVE_FILE_GROWTH ((0x00001000L))
value REG_FORCE_RESTORE ((0x00000008L))
value REG_FORCE_UNLOAD (1)
value REG_HIVE_EXACT_FILE_GROWTH ((0x00000080L))
value REG_HIVE_NO_RM ((0x00000100L))
value REG_HIVE_SINGLE_LOG ((0x00000200L))
value REG_IMMUTABLE ((0x00004000L))
value REG_LATEST_FORMAT (2)
value REG_LEGAL_CHANGE_FILTER ((REG_NOTIFY_CHANGE_NAME | REG_NOTIFY_CHANGE_ATTRIBUTES | REG_NOTIFY_CHANGE_LAST_SET | REG_NOTIFY_CHANGE_SECURITY | REG_NOTIFY_THREAD_AGNOSTIC))
value REG_LEGAL_OPTION ((REG_OPTION_RESERVED | REG_OPTION_NON_VOLATILE | REG_OPTION_VOLATILE | REG_OPTION_CREATE_LINK | REG_OPTION_BACKUP_RESTORE | REG_OPTION_OPEN_LINK | REG_OPTION_DONT_VIRTUALIZE))
value REG_LOAD_HIVE_OPEN_HANDLE ((0x00000800L))
value REG_MUI_STRING_TRUNCATE (0x00000001)
value REG_NOTIFY_CHANGE_ATTRIBUTES ((0x00000002L))
value REG_NOTIFY_CHANGE_LAST_SET ((0x00000004L))
value REG_NOTIFY_CHANGE_NAME ((0x00000001L))
value REG_NOTIFY_CHANGE_SECURITY ((0x00000008L))
value REG_NOTIFY_THREAD_AGNOSTIC ((0x10000000L))
value REG_NO_COMPRESSION (4)
value REG_NO_IMPERSONATION_FALLBACK ((0x00008000L))
value REG_NO_LAZY_FLUSH ((0x00000004L))
value REG_OPENED_EXISTING_KEY ((0x00000002L))
value REG_OPEN_LEGAL_OPTION ((REG_OPTION_RESERVED | REG_OPTION_BACKUP_RESTORE | REG_OPTION_OPEN_LINK | REG_OPTION_DONT_VIRTUALIZE))
value REG_OPEN_READ_ONLY ((0x00002000L))
value REG_OPTION_BACKUP_RESTORE ((0x00000004L))
value REG_OPTION_CREATE_LINK ((0x00000002L))
value REG_OPTION_DONT_VIRTUALIZE ((0x00000010L))
value REG_OPTION_NON_VOLATILE ((0x00000000L))
value REG_OPTION_OPEN_LINK ((0x00000008L))
value REG_OPTION_RESERVED ((0x00000000L))
value REG_OPTION_VOLATILE ((0x00000001L))
value REG_PROCESS_APPKEY (0x00000001)
value REG_PROCESS_PRIVATE ((0x00000020L))
value REG_REFRESH_HIVE ((0x00000002L))
value REG_SECURE_CONNECTION (1)
value REG_STANDARD_FORMAT (1)
value REG_START_JOURNAL ((0x00000040L))
value REG_UNLOAD_LEGAL_FLAGS ((REG_FORCE_UNLOAD))
value REG_USE_CURRENT_SECURITY_CONTEXT (0x00000002)
value REG_WHOLE_HIVE_VOLATILE ((0x00000001L))
value RELATIVE (2)
value REMOTE_NAME_INFO_LEVEL (0x00000002)
value REMOTE_PROTOCOL_INFO_FLAG_LOOPBACK (0x00000001)
value REMOTE_PROTOCOL_INFO_FLAG_OFFLINE (0x00000002)
value REMOTE_PROTOCOL_INFO_FLAG_PERSISTENT_HANDLE (0x00000004)
value REPLACEDLGORD (1541)
value REPLACEFILE_IGNORE_ACL_ERRORS (0x00000004)
value REPLACEFILE_IGNORE_MERGE_ERRORS (0x00000002)
value REPLACEFILE_WRITE_THROUGH (0x00000001)
value REPLACE_ALTERNATE (0xB)
value REPLACE_PRIMARY (0xA)
value REPORT_NOT_ABLE_TO_EXPORT_PRIVATE_KEY (0x0002)
value REPORT_NO_PRIVATE_KEY (0x0001)
value REQUEST_OPLOCK_CURRENT_VERSION (1)
value REQUEST_OPLOCK_INPUT_FLAG_ACK ((0x00000002))
value REQUEST_OPLOCK_INPUT_FLAG_COMPLETE_ACK_ON_CLOSE ((0x00000004))
value REQUEST_OPLOCK_INPUT_FLAG_REQUEST ((0x00000001))
value REQUEST_OPLOCK_OUTPUT_FLAG_ACK_REQUIRED ((0x00000001))
value REQUEST_OPLOCK_OUTPUT_FLAG_MODES_PROVIDED ((0x00000002))
value RESETDEV (7)
value RESOURCEDISPLAYTYPE_DIRECTORY (0x00000009)
value RESOURCEDISPLAYTYPE_DOMAIN (0x00000001)
value RESOURCEDISPLAYTYPE_FILE (0x00000004)
value RESOURCEDISPLAYTYPE_GENERIC (0x00000000)
value RESOURCEDISPLAYTYPE_GROUP (0x00000005)
value RESOURCEDISPLAYTYPE_NDSCONTAINER (0x0000000B)
value RESOURCEDISPLAYTYPE_NETWORK (0x00000006)
value RESOURCEDISPLAYTYPE_ROOT (0x00000007)
value RESOURCEDISPLAYTYPE_SERVER (0x00000002)
value RESOURCEDISPLAYTYPE_SHARE (0x00000003)
value RESOURCEDISPLAYTYPE_SHAREADMIN (0x00000008)
value RESOURCEDISPLAYTYPE_TREE (0x0000000A)
value RESOURCEMANAGER_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | RESOURCEMANAGER_GENERIC_READ | RESOURCEMANAGER_GENERIC_WRITE | RESOURCEMANAGER_GENERIC_EXECUTE))
value RESOURCEMANAGER_COMPLETE_PROPAGATION (( 0x0040 ))
value RESOURCEMANAGER_ENLIST (( 0x0008 ))
value RESOURCEMANAGER_GENERIC_EXECUTE ((STANDARD_RIGHTS_EXECUTE | RESOURCEMANAGER_RECOVER | RESOURCEMANAGER_ENLIST | RESOURCEMANAGER_GET_NOTIFICATION | RESOURCEMANAGER_COMPLETE_PROPAGATION | SYNCHRONIZE))
value RESOURCEMANAGER_GENERIC_READ ((STANDARD_RIGHTS_READ | RESOURCEMANAGER_QUERY_INFORMATION | SYNCHRONIZE))
value RESOURCEMANAGER_GENERIC_WRITE ((STANDARD_RIGHTS_WRITE | RESOURCEMANAGER_SET_INFORMATION | RESOURCEMANAGER_RECOVER | RESOURCEMANAGER_ENLIST | RESOURCEMANAGER_GET_NOTIFICATION | RESOURCEMANAGER_REGISTER_PROTOCOL | RESOURCEMANAGER_COMPLETE_PROPAGATION | SYNCHRONIZE))
value RESOURCEMANAGER_GET_NOTIFICATION (( 0x0010 ))
value RESOURCEMANAGER_QUERY_INFORMATION (( 0x0001 ))
value RESOURCEMANAGER_RECOVER (( 0x0004 ))
value RESOURCEMANAGER_REGISTER_PROTOCOL (( 0x0020 ))
value RESOURCEMANAGER_SET_INFORMATION (( 0x0002 ))
value RESOURCETYPE_ANY (0x00000000)
value RESOURCETYPE_DISK (0x00000001)
value RESOURCETYPE_PRINT (0x00000002)
value RESOURCETYPE_RESERVED (0x00000008)
value RESOURCETYPE_UNKNOWN (0xFFFFFFFF)
value RESOURCEUSAGE_ALL ((RESOURCEUSAGE_CONNECTABLE | RESOURCEUSAGE_CONTAINER | RESOURCEUSAGE_ATTACHED))
value RESOURCEUSAGE_ATTACHED (0x00000010)
value RESOURCEUSAGE_CONNECTABLE (0x00000001)
value RESOURCEUSAGE_CONTAINER (0x00000002)
value RESOURCEUSAGE_NOLOCALDEVICE (0x00000004)
value RESOURCEUSAGE_RESERVED (0x80000000)
value RESOURCEUSAGE_SIBLING (0x00000008)
value RESOURCE_CONNECTED (0x00000001)
value RESOURCE_CONTEXT (0x00000005)
value RESOURCE_ENUM_LN ((0x0001))
value RESOURCE_ENUM_MODULE_EXACT ((0x0010))
value RESOURCE_ENUM_MUI ((0x0002))
value RESOURCE_ENUM_MUI_SYSTEM ((0x0004))
value RESOURCE_ENUM_VALIDATE ((0x0008))
value RESOURCE_GLOBALNET (0x00000002)
value RESOURCE_MANAGER_COMMUNICATION (0x00000002)
value RESOURCE_MANAGER_MAXIMUM_OPTION (0x00000003)
value RESOURCE_MANAGER_VOLATILE (0x00000001)
value RESOURCE_RECENT (0x00000004)
value RESOURCE_REMEMBERED (0x00000003)
value RESTART_MAX_CMD_LINE (1024)
value RESTART_NO_CRASH (1)
value RESTART_NO_HANG (2)
value RESTART_NO_PATCH (4)
value RESTART_NO_REBOOT (8)
value RESTORE_CTM (4100)
value RESULT_IS_ADDED (0x0010)
value RESULT_IS_ALIAS (0x0001)
value RESULT_IS_CHANGED (0x0020)
value RESULT_IS_DELETED (0x0040)
value RES_CURSOR (2)
value RES_FLUSH_CACHE ((0x00000002))
value RES_ICON (1)
value RES_SERVICE ((0x00000004))
value RETRACT_IEPORT (3)
value RETURN_SMART_STATUS (0xDA)
value REVERSE_PRINT (( 0x00000001 ))
value REVISION_LENGTH (4)
value REVOCATION_OID_CRL_REVOCATION (((LPCSTR)1))
value RGB_GAMMA_MAX ((WORD)65000)
value RGB_GAMMA_MIN ((WORD)02500)
value RGN_AND (1)
value RGN_COPY (5)
value RGN_DIFF (4)
value RGN_ERROR (ERROR)
value RGN_MAX (RGN_COPY)
value RGN_MIN (RGN_AND)
value RGN_OR (2)
value RGN_XOR (3)
value RIDEV_APPKEYS (0x00000400)
value RIDEV_CAPTUREMOUSE (0x00000200)
value RIDEV_DEVNOTIFY (0x00002000)
value RIDEV_EXCLUDE (0x00000010)
value RIDEV_EXINPUTSINK (0x00001000)
value RIDEV_EXMODEMASK (0x000000F0)
value RIDEV_INPUTSINK (0x00000100)
value RIDEV_NOHOTKEYS (0x00000200)
value RIDEV_NOLEGACY (0x00000030)
value RIDEV_PAGEONLY (0x00000020)
value RIDEV_REMOVE (0x00000001)
value RIDI_DEVICEINFO (0x2000000b)
value RIDI_DEVICENAME (0x20000007)
value RIDI_PREPARSEDDATA (0x20000005)
value RID_HEADER (0x10000005)
value RID_INPUT (0x10000003)
value RIGHTMOST_BUTTON_PRESSED (0x0002)
value RIGHT_ALT_PRESSED (0x0001)
value RIGHT_CTRL_PRESSED (0x0004)
value RIM_INPUT (0)
value RIM_INPUTSINK (1)
value RIM_TYPEHID (2)
value RIM_TYPEKEYBOARD (1)
value RIM_TYPEMAX (2)
value RIM_TYPEMOUSE (0)
value RIP_EVENT (9)
value RI_KEY_BREAK (1)
value RI_KEY_MAKE (0)
value RI_KEY_TERMSRV_SET_LED (8)
value RI_KEY_TERMSRV_SHADOW (0x10)
value RI_MOUSE_HWHEEL (0x0800)
value RI_MOUSE_LEFT_BUTTON_DOWN (0x0001)
value RI_MOUSE_LEFT_BUTTON_UP (0x0002)
value RI_MOUSE_MIDDLE_BUTTON_DOWN (0x0010)
value RI_MOUSE_MIDDLE_BUTTON_UP (0x0020)
value RI_MOUSE_RIGHT_BUTTON_DOWN (0x0004)
value RI_MOUSE_RIGHT_BUTTON_UP (0x0008)
value RI_MOUSE_WHEEL (0x0400)
value ROTFLAGS_ALLOWANYCLIENT (0x2)
value ROTFLAGS_REGISTRATIONKEEPSALIVE (0x1)
value ROTREGFLAGS_ALLOWANYCLIENT (0x1)
value ROT_COMPARE_MAX (2048)
value RO_E_BLOCKED_CROSS_ASTA_CALL (_HRESULT_TYPEDEF_(0x8000001FL))
value RO_E_CANNOT_ACTIVATE_FULL_TRUST_SERVER (_HRESULT_TYPEDEF_(0x80000020L))
value RO_E_CANNOT_ACTIVATE_UNIVERSAL_APPLICATION_SERVER (_HRESULT_TYPEDEF_(0x80000021L))
value RO_E_CHANGE_NOTIFICATION_IN_PROGRESS (_HRESULT_TYPEDEF_(0x80000015L))
value RO_E_CLOSED (_HRESULT_TYPEDEF_(0x80000013L))
value RO_E_COMMITTED (_HRESULT_TYPEDEF_(0x8000001EL))
value RO_E_ERROR_STRING_NOT_FOUND (_HRESULT_TYPEDEF_(0x80000016L))
value RO_E_EXCLUSIVE_WRITE (_HRESULT_TYPEDEF_(0x80000014L))
value RO_E_INVALID_METADATA_FILE (_HRESULT_TYPEDEF_(0x80000012L))
value RO_E_METADATA_INVALID_TYPE_FORMAT (_HRESULT_TYPEDEF_(0x80000011L))
value RO_E_METADATA_NAME_IS_NAMESPACE (_HRESULT_TYPEDEF_(0x80000010L))
value RO_E_METADATA_NAME_NOT_FOUND (_HRESULT_TYPEDEF_(0x8000000FL))
value RO_E_MUST_BE_AGILE (_HRESULT_TYPEDEF_(0x8000001CL))
value RO_E_UNSUPPORTED_FROM_MTA (_HRESULT_TYPEDEF_(0x8000001DL))
value RPCFLG_ACCESS_LOCAL (0x00400000UL)
value RPCFLG_ASYNCHRONOUS (0x40000000UL)
value RPCFLG_AUTO_COMPLETE (0x08000000UL)
value RPCFLG_HAS_CALLBACK (0x04000000UL)
value RPCFLG_HAS_GUARANTEE (0x00000010UL)
value RPCFLG_HAS_MULTI_SYNTAXES (0x02000000UL)
value RPCFLG_INPUT_SYNCHRONOUS (0x20000000UL)
value RPCFLG_LOCAL_CALL (0x10000000UL)
value RPCFLG_MESSAGE (0x01000000UL)
value RPCFLG_NON_NDR (0x80000000UL)
value RPCFLG_SENDER_WAITING_FOR_REPLY (0x00800000UL)
value RPCFLG_WINRT_REMOTE_ASYNC (0x00000020UL)
value RPCNSAPI (DECLSPEC_IMPORT)
value RPCRTAPI (DECLSPEC_IMPORT)
value RPC_BHO_DONTLINGER ((0x2))
value RPC_BHO_EXCLUSIVE_AND_GUARANTEED ((0x4))
value RPC_BHO_NONCAUSAL ((0x1))
value RPC_BHT_OBJECT_UUID_VALID ((0x1))
value RPC_BUFFER_ASYNC (0x00008000)
value RPC_BUFFER_COMPLETE (0x00001000)
value RPC_BUFFER_EXTRA (0x00004000)
value RPC_BUFFER_NONOTIFY (0x00010000)
value RPC_BUFFER_PARTIAL (0x00002000)
value RPC_CALL_ATTRIBUTES_VERSION ((3))
value RPC_CALL_STATUS_CANCELLED (0x01)
value RPC_CALL_STATUS_DISCONNECTED (0x02)
value RPC_CONTEXT_HANDLE_DEFAULT_FLAGS (0x00000000UL)
value RPC_CONTEXT_HANDLE_DONT_SERIALIZE (0x20000000UL)
value RPC_CONTEXT_HANDLE_FLAGS (0x30000000UL)
value RPC_CONTEXT_HANDLE_SERIALIZE (0x10000000UL)
value RPC_C_AUTHN_CLOUD_AP (36)
value RPC_C_AUTHN_DCE_PRIVATE (1)
value RPC_C_AUTHN_DCE_PUBLIC (2)
value RPC_C_AUTHN_DEC_PUBLIC (4)
value RPC_C_AUTHN_DEFAULT (0xFFFFFFFFL)
value RPC_C_AUTHN_DIGEST (21)
value RPC_C_AUTHN_DPA (17)
value RPC_C_AUTHN_GSS_KERBEROS (16)
value RPC_C_AUTHN_GSS_NEGOTIATE (9)
value RPC_C_AUTHN_GSS_SCHANNEL (14)
value RPC_C_AUTHN_INFO_TYPE_HTTP (1)
value RPC_C_AUTHN_KERNEL (20)
value RPC_C_AUTHN_LEVEL_CALL (3)
value RPC_C_AUTHN_LEVEL_CONNECT (2)
value RPC_C_AUTHN_LEVEL_DEFAULT (0)
value RPC_C_AUTHN_LEVEL_NONE (1)
value RPC_C_AUTHN_LEVEL_PKT (4)
value RPC_C_AUTHN_LEVEL_PKT_INTEGRITY (5)
value RPC_C_AUTHN_LEVEL_PKT_PRIVACY (6)
value RPC_C_AUTHN_LIVEXP_SSP (35)
value RPC_C_AUTHN_LIVE_SSP (32)
value RPC_C_AUTHN_MQ (100)
value RPC_C_AUTHN_MSN (18)
value RPC_C_AUTHN_MSONLINE (82)
value RPC_C_AUTHN_NEGO_EXTENDER (30)
value RPC_C_AUTHN_NONE (0)
value RPC_C_AUTHN_WINNT (10)
value RPC_C_AUTHZ_DCE (2)
value RPC_C_AUTHZ_DEFAULT (0xffffffff)
value RPC_C_AUTHZ_NAME (1)
value RPC_C_AUTHZ_NONE (0)
value RPC_C_BINDING_DEFAULT_TIMEOUT (5)
value RPC_C_BINDING_INFINITE_TIMEOUT (10)
value RPC_C_BINDING_MAX_TIMEOUT (9)
value RPC_C_BINDING_MIN_TIMEOUT (0)
value RPC_C_BIND_TO_ALL_NICS (1)
value RPC_C_CANCEL_INFINITE_TIMEOUT (-1)
value RPC_C_DONT_FAIL (0x4)
value RPC_C_EP_ALL_ELTS (0)
value RPC_C_EP_MATCH_BY_BOTH (3)
value RPC_C_EP_MATCH_BY_IF (1)
value RPC_C_EP_MATCH_BY_OBJ (2)
value RPC_C_FULL_CERT_CHAIN (0x0001)
value RPC_C_HTTP_AUTHN_SCHEME_BASIC (0x00000001)
value RPC_C_HTTP_AUTHN_SCHEME_CERT (0x00010000)
value RPC_C_HTTP_AUTHN_SCHEME_DIGEST (0x00000008)
value RPC_C_HTTP_AUTHN_SCHEME_NEGOTIATE (0x00000010)
value RPC_C_HTTP_AUTHN_SCHEME_NTLM (0x00000002)
value RPC_C_HTTP_AUTHN_SCHEME_PASSPORT (0x00000004)
value RPC_C_HTTP_AUTHN_TARGET_PROXY (2)
value RPC_C_HTTP_AUTHN_TARGET_SERVER (1)
value RPC_C_HTTP_FLAG_ENABLE_CERT_REVOCATION_CHECK (16)
value RPC_C_HTTP_FLAG_IGNORE_CERT_CN_INVALID (8)
value RPC_C_HTTP_FLAG_USE_FIRST_AUTH_SCHEME (2)
value RPC_C_HTTP_FLAG_USE_SSL (1)
value RPC_C_IMP_LEVEL_ANONYMOUS (1)
value RPC_C_IMP_LEVEL_DEFAULT (0)
value RPC_C_IMP_LEVEL_DELEGATE (4)
value RPC_C_IMP_LEVEL_IDENTIFY (2)
value RPC_C_IMP_LEVEL_IMPERSONATE (3)
value RPC_C_INFINITE_TIMEOUT (INFINITE)
value RPC_C_LISTEN_MAX_CALLS_DEFAULT (1234)
value RPC_C_MGMT_INQ_IF_IDS (0)
value RPC_C_MGMT_INQ_PRINC_NAME (1)
value RPC_C_MGMT_INQ_STATS (2)
value RPC_C_MGMT_IS_SERVER_LISTEN (3)
value RPC_C_MGMT_STOP_SERVER_LISTEN (4)
value RPC_C_NOTIFY_ON_SEND_COMPLETE (0x1)
value RPC_C_NO_CREDENTIALS (((RPC_AUTH_IDENTITY_HANDLE) MAXUINT_PTR))
value RPC_C_NS_DEFAULT_EXP_AGE (-1)
value RPC_C_NS_SYNTAX_DCE (3)
value RPC_C_NS_SYNTAX_DEFAULT (0)
value RPC_C_OPT_ASYNC_BLOCK (15)
value RPC_C_OPT_BINDING_NONCAUSAL (9)
value RPC_C_OPT_CALL_TIMEOUT (12)
value RPC_C_OPT_COOKIE_AUTH ((7))
value RPC_C_OPT_DONT_LINGER (13)
value RPC_C_OPT_MAX_OPTIONS (17)
value RPC_C_OPT_OPTIMIZE_TIME (16)
value RPC_C_OPT_PRIVATE_BREAK_ON_SUSPEND (3)
value RPC_C_OPT_PRIVATE_DO_NOT_DISTURB (2)
value RPC_C_OPT_PRIVATE_SUPPRESS_WAKE (1)
value RPC_C_OPT_RESOURCE_TYPE_UUID ((8))
value RPC_C_OPT_SECURITY_CALLBACK (10)
value RPC_C_OPT_SESSION_ID ((6))
value RPC_C_OPT_TRANS_SEND_BUFFER_SIZE (5)
value RPC_C_OPT_TRUST_PEER (14)
value RPC_C_OPT_UNIQUE_BINDING (11)
value RPC_C_PARM_BUFFER_LENGTH (2)
value RPC_C_PARM_MAX_PACKET_LENGTH (1)
value RPC_C_PROFILE_ALL_ELT (1)
value RPC_C_PROFILE_ALL_ELTS (RPC_C_PROFILE_ALL_ELT)
value RPC_C_PROFILE_DEFAULT_ELT (0)
value RPC_C_PROFILE_MATCH_BY_BOTH (4)
value RPC_C_PROFILE_MATCH_BY_IF (2)
value RPC_C_PROFILE_MATCH_BY_MBR (3)
value RPC_C_PROTECT_LEVEL_CALL ((RPC_C_AUTHN_LEVEL_CALL))
value RPC_C_PROTECT_LEVEL_CONNECT ((RPC_C_AUTHN_LEVEL_CONNECT))
value RPC_C_PROTECT_LEVEL_DEFAULT ((RPC_C_AUTHN_LEVEL_DEFAULT))
value RPC_C_PROTECT_LEVEL_NONE ((RPC_C_AUTHN_LEVEL_NONE))
value RPC_C_PROTECT_LEVEL_PKT ((RPC_C_AUTHN_LEVEL_PKT))
value RPC_C_PROTECT_LEVEL_PKT_INTEGRITY ((RPC_C_AUTHN_LEVEL_PKT_INTEGRITY))
value RPC_C_PROTECT_LEVEL_PKT_PRIVACY ((RPC_C_AUTHN_LEVEL_PKT_PRIVACY))
value RPC_C_PROTSEQ_MAX_REQS_DEFAULT (10)
value RPC_C_QOS_CAPABILITIES_ANY_AUTHORITY (0x4)
value RPC_C_QOS_CAPABILITIES_DEFAULT (0x0)
value RPC_C_QOS_CAPABILITIES_IGNORE_DELEGATE_FAILURE (0x8)
value RPC_C_QOS_CAPABILITIES_LOCAL_MA_HINT (0x10)
value RPC_C_QOS_CAPABILITIES_MAKE_FULLSIC (0x2)
value RPC_C_QOS_CAPABILITIES_MUTUAL_AUTH (0x1)
value RPC_C_QOS_CAPABILITIES_SCHANNEL_FULL_AUTH_IDENTITY (0x20)
value RPC_C_QOS_IDENTITY_DYNAMIC (1)
value RPC_C_QOS_IDENTITY_STATIC (0)
value RPC_C_RPCHTTP_USE_LOAD_BALANCE (0x8)
value RPC_C_SECURITY_QOS_VERSION (1)
value RPC_C_STATS_CALLS_IN (0)
value RPC_C_STATS_CALLS_OUT (1)
value RPC_C_STATS_PKTS_IN (2)
value RPC_C_STATS_PKTS_OUT (3)
value RPC_C_TRY_ENFORCE_MAX_CALLS (0x10)
value RPC_C_USE_INTERNET_PORT (0x1)
value RPC_C_USE_INTRANET_PORT (0x2)
value RPC_C_VERS_ALL (1)
value RPC_C_VERS_COMPATIBLE (2)
value RPC_C_VERS_EXACT (3)
value RPC_C_VERS_MAJOR_ONLY (4)
value RPC_C_VERS_UPTO (5)
value RPC_EEINFO_VERSION (1)
value RPC_ENDPOINT_TEMPLATE (RPC_ENDPOINT_TEMPLATEA)
value RPC_E_ACCESS_DENIED (_HRESULT_TYPEDEF_(0x8001011BL))
value RPC_E_ATTEMPTED_MULTITHREAD (_HRESULT_TYPEDEF_(0x80010102L))
value RPC_E_CALL_CANCELED (_HRESULT_TYPEDEF_(0x80010002L))
value RPC_E_CALL_COMPLETE (_HRESULT_TYPEDEF_(0x80010117L))
value RPC_E_CALL_REJECTED (_HRESULT_TYPEDEF_(0x80010001L))
value RPC_E_CANTCALLOUT_AGAIN (_HRESULT_TYPEDEF_(0x80010011L))
value RPC_E_CANTCALLOUT_INASYNCCALL (_HRESULT_TYPEDEF_(0x80010004L))
value RPC_E_CANTCALLOUT_INEXTERNALCALL (_HRESULT_TYPEDEF_(0x80010005L))
value RPC_E_CANTCALLOUT_ININPUTSYNCCALL (_HRESULT_TYPEDEF_(0x8001010DL))
value RPC_E_CANTPOST_INSENDCALL (_HRESULT_TYPEDEF_(0x80010003L))
value RPC_E_CANTTRANSMIT_CALL (_HRESULT_TYPEDEF_(0x8001000AL))
value RPC_E_CHANGED_MODE (_HRESULT_TYPEDEF_(0x80010106L))
value RPC_E_CLIENT_CANTMARSHAL_DATA (_HRESULT_TYPEDEF_(0x8001000BL))
value RPC_E_CLIENT_CANTUNMARSHAL_DATA (_HRESULT_TYPEDEF_(0x8001000CL))
value RPC_E_CLIENT_DIED (_HRESULT_TYPEDEF_(0x80010008L))
value RPC_E_CONNECTION_TERMINATED (_HRESULT_TYPEDEF_(0x80010006L))
value RPC_E_DISCONNECTED (_HRESULT_TYPEDEF_(0x80010108L))
value RPC_E_FAULT (_HRESULT_TYPEDEF_(0x80010104L))
value RPC_E_FULLSIC_REQUIRED (_HRESULT_TYPEDEF_(0x80010121L))
value RPC_E_INVALIDMETHOD (_HRESULT_TYPEDEF_(0x80010107L))
value RPC_E_INVALID_CALLDATA (_HRESULT_TYPEDEF_(0x8001010CL))
value RPC_E_INVALID_DATA (_HRESULT_TYPEDEF_(0x8001000FL))
value RPC_E_INVALID_DATAPACKET (_HRESULT_TYPEDEF_(0x80010009L))
value RPC_E_INVALID_EXTENSION (_HRESULT_TYPEDEF_(0x80010112L))
value RPC_E_INVALID_HEADER (_HRESULT_TYPEDEF_(0x80010111L))
value RPC_E_INVALID_IPID (_HRESULT_TYPEDEF_(0x80010113L))
value RPC_E_INVALID_OBJECT (_HRESULT_TYPEDEF_(0x80010114L))
value RPC_E_INVALID_OBJREF (_HRESULT_TYPEDEF_(0x8001011DL))
value RPC_E_INVALID_PARAMETER (_HRESULT_TYPEDEF_(0x80010010L))
value RPC_E_INVALID_STD_NAME (_HRESULT_TYPEDEF_(0x80010122L))
value RPC_E_NOT_REGISTERED (_HRESULT_TYPEDEF_(0x80010103L))
value RPC_E_NO_CONTEXT (_HRESULT_TYPEDEF_(0x8001011EL))
value RPC_E_NO_GOOD_SECURITY_PACKAGES (_HRESULT_TYPEDEF_(0x8001011AL))
value RPC_E_NO_SYNC (_HRESULT_TYPEDEF_(0x80010120L))
value RPC_E_OUT_OF_RESOURCES (_HRESULT_TYPEDEF_(0x80010101L))
value RPC_E_REMOTE_DISABLED (_HRESULT_TYPEDEF_(0x8001011CL))
value RPC_E_RETRY (_HRESULT_TYPEDEF_(0x80010109L))
value RPC_E_SERVERCALL_REJECTED (_HRESULT_TYPEDEF_(0x8001010BL))
value RPC_E_SERVERCALL_RETRYLATER (_HRESULT_TYPEDEF_(0x8001010AL))
value RPC_E_SERVERFAULT (_HRESULT_TYPEDEF_(0x80010105L))
value RPC_E_SERVER_CANTMARSHAL_DATA (_HRESULT_TYPEDEF_(0x8001000DL))
value RPC_E_SERVER_CANTUNMARSHAL_DATA (_HRESULT_TYPEDEF_(0x8001000EL))
value RPC_E_SERVER_DIED (_HRESULT_TYPEDEF_(0x80010007L))
value RPC_E_SERVER_DIED_DNE (_HRESULT_TYPEDEF_(0x80010012L))
value RPC_E_SYS_CALL_FAILED (_HRESULT_TYPEDEF_(0x80010100L))
value RPC_E_THREAD_NOT_INIT (_HRESULT_TYPEDEF_(0x8001010FL))
value RPC_E_TIMEOUT (_HRESULT_TYPEDEF_(0x8001011FL))
value RPC_E_TOO_LATE (_HRESULT_TYPEDEF_(0x80010119L))
value RPC_E_UNEXPECTED (_HRESULT_TYPEDEF_(0x8001FFFFL))
value RPC_E_UNSECURE_CALL (_HRESULT_TYPEDEF_(0x80010118L))
value RPC_E_VERSION_MISMATCH (_HRESULT_TYPEDEF_(0x80010110L))
value RPC_E_WRONG_THREAD (_HRESULT_TYPEDEF_(0x8001010EL))
value RPC_FLAGS_VALID_BIT (0x00008000)
value RPC_FW_IF_FLAG_DCOM (0x0001)
value RPC_HTTP_TRANSPORT_CREDENTIALS (RPC_HTTP_TRANSPORT_CREDENTIALS_A)
value RPC_IF_ALLOW_CALLBACKS_WITH_NO_AUTH (0x0010)
value RPC_IF_ALLOW_LOCAL_ONLY (0x0020)
value RPC_IF_ALLOW_SECURE_ONLY (0x0008)
value RPC_IF_ALLOW_UNKNOWN_AUTHORITY (0x0004)
value RPC_IF_ASYNC_CALLBACK (0x0100)
value RPC_IF_AUTOLISTEN (0x0001)
value RPC_IF_OLE (0x0002)
value RPC_IF_SEC_CACHE_PER_PROC (0x0080)
value RPC_IF_SEC_NO_CACHE (0x0040)
value RPC_INTERFACE_HAS_PIPES (0x0001)
value RPC_INTERFACE_TEMPLATE (RPC_INTERFACE_TEMPLATEA)
value RPC_NCA_FLAGS_BROADCAST (0x00000002)
value RPC_NCA_FLAGS_DEFAULT (0x00000000)
value RPC_NCA_FLAGS_IDEMPOTENT (0x00000001)
value RPC_NCA_FLAGS_MAYBE (0x00000004)
value RPC_PROTSEQ_HTTP ((0x4))
value RPC_PROTSEQ_LRPC ((0x3))
value RPC_PROTSEQ_NMP ((0x2))
value RPC_PROTSEQ_TCP ((0x1))
value RPC_PROTSEQ_VECTOR (RPC_PROTSEQ_VECTORA)
value RPC_PROXY_CONNECTION_TYPE_IN_PROXY (0)
value RPC_PROXY_CONNECTION_TYPE_OUT_PROXY (1)
value RPC_QUERY_CALL_LOCAL_ADDRESS ((0x08))
value RPC_QUERY_CLIENT_ID ((0x80))
value RPC_QUERY_CLIENT_PID ((0x10))
value RPC_QUERY_CLIENT_PRINCIPAL_NAME ((0x04))
value RPC_QUERY_IS_CLIENT_LOCAL ((0x20))
value RPC_QUERY_NO_AUTH_REQUIRED ((0x40))
value RPC_QUERY_SERVER_PRINCIPAL_NAME ((0x02))
value RPC_SYSTEM_HANDLE_FREE_ALL (3)
value RPC_SYSTEM_HANDLE_FREE_ERROR_ON_CLOSE (4)
value RPC_SYSTEM_HANDLE_FREE_RETRIEVED (2)
value RPC_SYSTEM_HANDLE_FREE_UNRETRIEVED (1)
value RPC_S_ACCESS_DENIED (ERROR_ACCESS_DENIED)
value RPC_S_ADDRESS_ERROR (1768)
value RPC_S_ALREADY_LISTENING (1713)
value RPC_S_ALREADY_REGISTERED (1711)
value RPC_S_ASYNC_CALL_PENDING (ERROR_IO_PENDING)
value RPC_S_BINDING_HAS_NO_AUTH (1746)
value RPC_S_BINDING_INCOMPLETE (1819)
value RPC_S_BUFFER_TOO_SMALL (ERROR_INSUFFICIENT_BUFFER)
value RPC_S_CALLPENDING (_HRESULT_TYPEDEF_(0x80010115L))
value RPC_S_CALL_CANCELLED (1818)
value RPC_S_CALL_FAILED (1726)
value RPC_S_CALL_FAILED_DNE (1727)
value RPC_S_CALL_IN_PROGRESS (1791)
value RPC_S_CANNOT_SUPPORT (1764)
value RPC_S_CANT_CREATE_ENDPOINT (1720)
value RPC_S_COMM_FAILURE (1820)
value RPC_S_COOKIE_AUTH_FAILED (1833)
value RPC_S_DO_NOT_DISTURB (1834)
value RPC_S_DUPLICATE_ENDPOINT (1740)
value RPC_S_ENTRY_ALREADY_EXISTS (1760)
value RPC_S_ENTRY_NOT_FOUND (1761)
value RPC_S_ENTRY_TYPE_MISMATCH (1922)
value RPC_S_FP_DIV_ZERO (1769)
value RPC_S_FP_OVERFLOW (1771)
value RPC_S_FP_UNDERFLOW (1770)
value RPC_S_GROUP_MEMBER_NOT_FOUND (1898)
value RPC_S_GRP_ELT_NOT_ADDED (1928)
value RPC_S_GRP_ELT_NOT_REMOVED (1929)
value RPC_S_INCOMPLETE_NAME (1755)
value RPC_S_INTERFACE_NOT_EXPORTED (1924)
value RPC_S_INTERFACE_NOT_FOUND (1759)
value RPC_S_INTERNAL_ERROR (1766)
value RPC_S_INVALID_ARG (ERROR_INVALID_PARAMETER)
value RPC_S_INVALID_ASYNC_CALL (1915)
value RPC_S_INVALID_ASYNC_HANDLE (1914)
value RPC_S_INVALID_AUTH_IDENTITY (1749)
value RPC_S_INVALID_BINDING (1702)
value RPC_S_INVALID_BOUND (1734)
value RPC_S_INVALID_ENDPOINT_FORMAT (1706)
value RPC_S_INVALID_LEVEL (ERROR_INVALID_PARAMETER)
value RPC_S_INVALID_NAF_ID (1763)
value RPC_S_INVALID_NAME_SYNTAX (1736)
value RPC_S_INVALID_NETWORK_OPTIONS (1724)
value RPC_S_INVALID_NET_ADDR (1707)
value RPC_S_INVALID_OBJECT (1900)
value RPC_S_INVALID_RPC_PROTSEQ (1704)
value RPC_S_INVALID_SECURITY_DESC (ERROR_INVALID_SECURITY_DESCR)
value RPC_S_INVALID_STRING_BINDING (1700)
value RPC_S_INVALID_STRING_UUID (1705)
value RPC_S_INVALID_TAG (1733)
value RPC_S_INVALID_TIMEOUT (1709)
value RPC_S_INVALID_VERS_OPTION (1756)
value RPC_S_MAX_CALLS_TOO_SMALL (1742)
value RPC_S_NAME_SERVICE_UNAVAILABLE (1762)
value RPC_S_NOTHING_TO_EXPORT (1754)
value RPC_S_NOT_ALL_OBJS_EXPORTED (1923)
value RPC_S_NOT_ALL_OBJS_UNEXPORTED (1758)
value RPC_S_NOT_CANCELLED (1826)
value RPC_S_NOT_ENOUGH_QUOTA (ERROR_NOT_ENOUGH_QUOTA)
value RPC_S_NOT_LISTENING (1715)
value RPC_S_NOT_RPC_ERROR (1823)
value RPC_S_NO_BINDINGS (1718)
value RPC_S_NO_CALL_ACTIVE (1725)
value RPC_S_NO_CONTEXT_AVAILABLE (1765)
value RPC_S_NO_ENDPOINT_FOUND (1708)
value RPC_S_NO_ENTRY_NAME (1735)
value RPC_S_NO_INTERFACES (1817)
value RPC_S_NO_MORE_BINDINGS (1806)
value RPC_S_NO_MORE_MEMBERS (1757)
value RPC_S_NO_PRINC_NAME (1822)
value RPC_S_NO_PROTSEQS (1719)
value RPC_S_NO_PROTSEQS_REGISTERED (1714)
value RPC_S_OBJECT_NOT_FOUND (1710)
value RPC_S_OK (ERROR_SUCCESS)
value RPC_S_OUT_OF_MEMORY (ERROR_OUTOFMEMORY)
value RPC_S_OUT_OF_RESOURCES (1721)
value RPC_S_OUT_OF_THREADS (ERROR_MAX_THRDS_REACHED)
value RPC_S_PRF_ELT_NOT_ADDED (1926)
value RPC_S_PRF_ELT_NOT_REMOVED (1927)
value RPC_S_PROCNUM_OUT_OF_RANGE (1745)
value RPC_S_PROFILE_NOT_ADDED (1925)
value RPC_S_PROTOCOL_ERROR (1728)
value RPC_S_PROTSEQ_NOT_FOUND (1744)
value RPC_S_PROTSEQ_NOT_SUPPORTED (1703)
value RPC_S_PROXY_ACCESS_DENIED (1729)
value RPC_S_RUNTIME_UNINITIALIZED (ERROR_INVALID_FUNCTION)
value RPC_S_SEC_PKG_ERROR (1825)
value RPC_S_SEND_INCOMPLETE (1913)
value RPC_S_SERVER_OUT_OF_MEMORY (ERROR_NOT_ENOUGH_SERVER_MEMORY)
value RPC_S_SERVER_TOO_BUSY (1723)
value RPC_S_SERVER_UNAVAILABLE (1722)
value RPC_S_STRING_TOO_LONG (1743)
value RPC_S_SYSTEM_HANDLE_COUNT_EXCEEDED (1835)
value RPC_S_SYSTEM_HANDLE_TYPE_MISMATCH (1836)
value RPC_S_TIMEOUT (ERROR_TIMEOUT)
value RPC_S_TYPE_ALREADY_REGISTERED (1712)
value RPC_S_UNKNOWN_AUTHN_LEVEL (1748)
value RPC_S_UNKNOWN_AUTHN_SERVICE (1747)
value RPC_S_UNKNOWN_AUTHN_TYPE (1741)
value RPC_S_UNKNOWN_AUTHZ_SERVICE (1750)
value RPC_S_UNKNOWN_IF (1717)
value RPC_S_UNKNOWN_MGR_TYPE (1716)
value RPC_S_UNKNOWN_PRINCIPAL (ERROR_NONE_MAPPED)
value RPC_S_UNSUPPORTED_AUTHN_LEVEL (1821)
value RPC_S_UNSUPPORTED_NAME_SYNTAX (1737)
value RPC_S_UNSUPPORTED_TRANS_SYN (1730)
value RPC_S_UNSUPPORTED_TYPE (1732)
value RPC_S_UUID_LOCAL_ONLY (1824)
value RPC_S_UUID_NO_ADDRESS (1739)
value RPC_S_WAITONTIMER (_HRESULT_TYPEDEF_(0x80010116L))
value RPC_S_WRONG_KIND_OF_BINDING (1701)
value RPC_S_ZERO_DIVIDE (1767)
value RPC_TYPE_DISCONNECT_EVENT_CONTEXT_HANDLE (0x80000000UL)
value RPC_TYPE_STRICT_CONTEXT_HANDLE (0x40000000UL)
value RPC_X_BAD_STUB_DATA (1783)
value RPC_X_BYTE_COUNT_TOO_SMALL (1782)
value RPC_X_ENUM_VALUE_OUT_OF_RANGE (1781)
value RPC_X_ENUM_VALUE_TOO_LARGE (RPC_X_ENUM_VALUE_OUT_OF_RANGE)
value RPC_X_INVALID_BOUND (RPC_S_INVALID_BOUND)
value RPC_X_INVALID_BUFFER (ERROR_INVALID_USER_BUFFER)
value RPC_X_INVALID_ES_ACTION (1827)
value RPC_X_INVALID_PIPE_OBJECT (1830)
value RPC_X_INVALID_PIPE_OPERATION (RPC_X_WRONG_PIPE_ORDER)
value RPC_X_INVALID_TAG (RPC_S_INVALID_TAG)
value RPC_X_NO_MEMORY (RPC_S_OUT_OF_MEMORY)
value RPC_X_NO_MORE_ENTRIES (1772)
value RPC_X_NULL_REF_POINTER (1780)
value RPC_X_PIPE_APP_MEMORY (ERROR_OUTOFMEMORY)
value RPC_X_PIPE_CLOSED (1916)
value RPC_X_PIPE_DISCIPLINE_ERROR (1917)
value RPC_X_PIPE_EMPTY (1918)
value RPC_X_SS_CANNOT_GET_CALL_HANDLE (1779)
value RPC_X_SS_CHAR_TRANS_OPEN_FAIL (1773)
value RPC_X_SS_CHAR_TRANS_SHORT_FILE (1774)
value RPC_X_SS_CONTEXT_DAMAGED (1777)
value RPC_X_SS_CONTEXT_MISMATCH (ERROR_INVALID_HANDLE)
value RPC_X_SS_HANDLES_MISMATCH (1778)
value RPC_X_SS_IN_NULL_CONTEXT (1775)
value RPC_X_WRONG_ES_VERSION (1828)
value RPC_X_WRONG_PIPE_ORDER (1831)
value RPC_X_WRONG_PIPE_VERSION (1832)
value RPC_X_WRONG_STUB_VERSION (1829)
value RRF_NOEXPAND (0x10000000)
value RRF_RT_ANY (0x0000ffff)
value RRF_RT_DWORD ((RRF_RT_REG_BINARY | RRF_RT_REG_DWORD))
value RRF_RT_QWORD ((RRF_RT_REG_BINARY | RRF_RT_REG_QWORD))
value RRF_RT_REG_BINARY (0x00000008)
value RRF_RT_REG_DWORD (0x00000010)
value RRF_RT_REG_EXPAND_SZ (0x00000004)
value RRF_RT_REG_MULTI_SZ (0x00000020)
value RRF_RT_REG_NONE (0x00000001)
value RRF_RT_REG_QWORD (0x00000040)
value RRF_RT_REG_SZ (0x00000002)
value RRF_ZEROONFAILURE (0x20000000)
value RSA_CSP_PUBLICKEYBLOB (((LPCSTR) 19))
value RTL_CONDITION_VARIABLE_LOCKMODE_SHARED (0x1)
value RTL_CORRELATION_VECTOR_STRING_LENGTH (129)
value RTL_CORRELATION_VECTOR_VERSION_CURRENT (RTL_CORRELATION_VECTOR_VERSION_2)
value RTL_CRITICAL_SECTION_ALL_FLAG_BITS (0xFF000000)
value RTL_CRITICAL_SECTION_DEBUG_FLAG_STATIC_INIT (0x00000001)
value RTL_CRITICAL_SECTION_FLAG_DYNAMIC_SPIN (0x02000000)
value RTL_CRITICAL_SECTION_FLAG_FORCE_DEBUG_INFO (0x10000000)
value RTL_CRITICAL_SECTION_FLAG_NO_DEBUG_INFO (0x01000000)
value RTL_CRITICAL_SECTION_FLAG_RESOURCE_TYPE (0x08000000)
value RTL_CRITICAL_SECTION_FLAG_STATIC_INIT (0x04000000)
value RTL_RUN_ONCE_ASYNC (0x00000002UL)
value RTL_RUN_ONCE_CHECK_ONLY (0x00000001UL)
value RTL_RUN_ONCE_CTX_RESERVED_BITS (2)
value RTL_RUN_ONCE_INIT_FAILED (0x00000004UL)
value RTL_UMS_VERSION ((0x0100))
value RTS_CONTROL_DISABLE (0x00)
value RTS_CONTROL_ENABLE (0x01)
value RTS_CONTROL_HANDSHAKE (0x02)
value RTS_CONTROL_TOGGLE (0x03)
value RT_ACCELERATOR (MAKEINTRESOURCE(9))
value RT_ANICURSOR (MAKEINTRESOURCE(21))
value RT_ANIICON (MAKEINTRESOURCE(22))
value RT_BITMAP (MAKEINTRESOURCE(2))
value RT_CURSOR (MAKEINTRESOURCE(1))
value RT_DIALOG (MAKEINTRESOURCE(5))
value RT_DLGINCLUDE (MAKEINTRESOURCE(17))
value RT_FONT (MAKEINTRESOURCE(8))
value RT_FONTDIR (MAKEINTRESOURCE(7))
value RT_GROUP_CURSOR (MAKEINTRESOURCE((ULONG_PTR)(RT_CURSOR) + DIFFERENCE))
value RT_GROUP_ICON (MAKEINTRESOURCE((ULONG_PTR)(RT_ICON) + DIFFERENCE))
value RT_HTML (MAKEINTRESOURCE(23))
value RT_ICON (MAKEINTRESOURCE(3))
value RT_MANIFEST (MAKEINTRESOURCE(24))
value RT_MENU (MAKEINTRESOURCE(4))
value RT_MESSAGETABLE (MAKEINTRESOURCE(11))
value RT_PLUGPLAY (MAKEINTRESOURCE(19))
value RT_RCDATA (MAKEINTRESOURCE(10))
value RT_STRING (MAKEINTRESOURCE(6))
value RT_VERSION (MAKEINTRESOURCE(16))
value RT_VXD (MAKEINTRESOURCE(20))
value RUNDLGORD (1545)
value RUNTIME_FUNCTION_INDIRECT (0x1)
value RUSSIAN_CHARSET (204)
value SACL_SECURITY_INFORMATION ((0x00000008L))
value SANDBOX_INERT (0x2)
value SAVE_ATTRIBUTE_VALUES (0xD3)
value SAVE_CTM (4101)
value SBM_ENABLE_ARROWS (0x00E4)
value SBM_GETPOS (0x00E1)
value SBM_GETRANGE (0x00E3)
value SBM_GETSCROLLBARINFO (0x00EB)
value SBM_GETSCROLLINFO (0x00EA)
value SBM_SETPOS (0x00E0)
value SBM_SETRANGE (0x00E2)
value SBM_SETRANGEREDRAW (0x00E6)
value SBM_SETSCROLLINFO (0x00E9)
value SBS_BOTTOMALIGN (0x0004L)
value SBS_HORZ (0x0000L)
value SBS_LEFTALIGN (0x0002L)
value SBS_RIGHTALIGN (0x0004L)
value SBS_SIZEBOX (0x0008L)
value SBS_SIZEBOXBOTTOMRIGHTALIGN (0x0004L)
value SBS_SIZEBOXTOPLEFTALIGN (0x0002L)
value SBS_SIZEGRIP (0x0010L)
value SBS_TOPALIGN (0x0002L)
value SBS_VERT (0x0001L)
value SB_BOTH (3)
value SB_BOTTOM (7)
value SB_CONST_ALPHA (0x00000001)
value SB_CTL (2)
value SB_ENDSCROLL (8)
value SB_GRAD_RECT (0x00000010)
value SB_GRAD_TRI (0x00000020)
value SB_HORZ (0)
value SB_LEFT (6)
value SB_LINEDOWN (1)
value SB_LINELEFT (0)
value SB_LINERIGHT (1)
value SB_LINEUP (0)
value SB_NONE (0x00000000)
value SB_PAGEDOWN (3)
value SB_PAGELEFT (2)
value SB_PAGERIGHT (3)
value SB_PAGEUP (2)
value SB_PIXEL_ALPHA (0x00000002)
value SB_PREMULT_ALPHA (0x00000004)
value SB_RIGHT (7)
value SB_THUMBPOSITION (4)
value SB_THUMBTRACK (5)
value SB_TOP (6)
value SB_VERT (1)
value SCALINGFACTORX (114)
value SCALINGFACTORY (115)
value SCARD_ABSENT (1)
value SCARD_ATR_LENGTH (33)
value SCARD_ATTR_DEVICE_FRIENDLY_NAME (SCARD_ATTR_DEVICE_FRIENDLY_NAME_A)
value SCARD_ATTR_DEVICE_SYSTEM_NAME (SCARD_ATTR_DEVICE_SYSTEM_NAME_A)
value SCARD_AUDIT_CHV_FAILURE (0x0)
value SCARD_AUDIT_CHV_SUCCESS (0x1)
value SCARD_AUTOALLOCATE ((DWORD)(-1))
value SCARD_CLASS_COMMUNICATIONS (2)
value SCARD_CLASS_ICC_STATE (9)
value SCARD_CLASS_IFD_PROTOCOL (8)
value SCARD_CLASS_MECHANICAL (6)
value SCARD_CLASS_PERF (0x7ffe)
value SCARD_CLASS_POWER_MGMT (4)
value SCARD_CLASS_PROTOCOL (3)
value SCARD_CLASS_SECURITY (5)
value SCARD_CLASS_SYSTEM (0x7fff)
value SCARD_CLASS_VENDOR_DEFINED (7)
value SCARD_CLASS_VENDOR_INFO (1)
value SCARD_COLD_RESET (1)
value SCARD_EJECT_CARD (3)
value SCARD_E_BAD_SEEK (_HRESULT_TYPEDEF_(0x80100029L))
value SCARD_E_CANCELLED (_HRESULT_TYPEDEF_(0x80100002L))
value SCARD_E_CANT_DISPOSE (_HRESULT_TYPEDEF_(0x8010000EL))
value SCARD_E_CARD_UNSUPPORTED (_HRESULT_TYPEDEF_(0x8010001CL))
value SCARD_E_CERTIFICATE_UNAVAILABLE (_HRESULT_TYPEDEF_(0x8010002DL))
value SCARD_E_COMM_DATA_LOST (_HRESULT_TYPEDEF_(0x8010002FL))
value SCARD_E_DIR_NOT_FOUND (_HRESULT_TYPEDEF_(0x80100023L))
value SCARD_E_DUPLICATE_READER (_HRESULT_TYPEDEF_(0x8010001BL))
value SCARD_E_FILE_NOT_FOUND (_HRESULT_TYPEDEF_(0x80100024L))
value SCARD_E_ICC_CREATEORDER (_HRESULT_TYPEDEF_(0x80100021L))
value SCARD_E_ICC_INSTALLATION (_HRESULT_TYPEDEF_(0x80100020L))
value SCARD_E_INSUFFICIENT_BUFFER (_HRESULT_TYPEDEF_(0x80100008L))
value SCARD_E_INVALID_ATR (_HRESULT_TYPEDEF_(0x80100015L))
value SCARD_E_INVALID_CHV (_HRESULT_TYPEDEF_(0x8010002AL))
value SCARD_E_INVALID_HANDLE (_HRESULT_TYPEDEF_(0x80100003L))
value SCARD_E_INVALID_PARAMETER (_HRESULT_TYPEDEF_(0x80100004L))
value SCARD_E_INVALID_TARGET (_HRESULT_TYPEDEF_(0x80100005L))
value SCARD_E_INVALID_VALUE (_HRESULT_TYPEDEF_(0x80100011L))
value SCARD_E_NOT_READY (_HRESULT_TYPEDEF_(0x80100010L))
value SCARD_E_NOT_TRANSACTED (_HRESULT_TYPEDEF_(0x80100016L))
value SCARD_E_NO_ACCESS (_HRESULT_TYPEDEF_(0x80100027L))
value SCARD_E_NO_DIR (_HRESULT_TYPEDEF_(0x80100025L))
value SCARD_E_NO_FILE (_HRESULT_TYPEDEF_(0x80100026L))
value SCARD_E_NO_KEY_CONTAINER (_HRESULT_TYPEDEF_(0x80100030L))
value SCARD_E_NO_MEMORY (_HRESULT_TYPEDEF_(0x80100006L))
value SCARD_E_NO_PIN_CACHE (_HRESULT_TYPEDEF_(0x80100033L))
value SCARD_E_NO_READERS_AVAILABLE (_HRESULT_TYPEDEF_(0x8010002EL))
value SCARD_E_NO_SERVICE (_HRESULT_TYPEDEF_(0x8010001DL))
value SCARD_E_NO_SMARTCARD (_HRESULT_TYPEDEF_(0x8010000CL))
value SCARD_E_NO_SUCH_CERTIFICATE (_HRESULT_TYPEDEF_(0x8010002CL))
value SCARD_E_PCI_TOO_SMALL (_HRESULT_TYPEDEF_(0x80100019L))
value SCARD_E_PIN_CACHE_EXPIRED (_HRESULT_TYPEDEF_(0x80100032L))
value SCARD_E_PROTO_MISMATCH (_HRESULT_TYPEDEF_(0x8010000FL))
value SCARD_E_READER_UNAVAILABLE (_HRESULT_TYPEDEF_(0x80100017L))
value SCARD_E_READER_UNSUPPORTED (_HRESULT_TYPEDEF_(0x8010001AL))
value SCARD_E_READ_ONLY_CARD (_HRESULT_TYPEDEF_(0x80100034L))
value SCARD_E_SERVER_TOO_BUSY (_HRESULT_TYPEDEF_(0x80100031L))
value SCARD_E_SERVICE_STOPPED (_HRESULT_TYPEDEF_(0x8010001EL))
value SCARD_E_SHARING_VIOLATION (_HRESULT_TYPEDEF_(0x8010000BL))
value SCARD_E_SYSTEM_CANCELLED (_HRESULT_TYPEDEF_(0x80100012L))
value SCARD_E_TIMEOUT (_HRESULT_TYPEDEF_(0x8010000AL))
value SCARD_E_UNEXPECTED (_HRESULT_TYPEDEF_(0x8010001FL))
value SCARD_E_UNKNOWN_CARD (_HRESULT_TYPEDEF_(0x8010000DL))
value SCARD_E_UNKNOWN_READER (_HRESULT_TYPEDEF_(0x80100009L))
value SCARD_E_UNKNOWN_RES_MNG (_HRESULT_TYPEDEF_(0x8010002BL))
value SCARD_E_UNSUPPORTED_FEATURE (_HRESULT_TYPEDEF_(0x80100022L))
value SCARD_E_WRITE_TOO_MANY (_HRESULT_TYPEDEF_(0x80100028L))
value SCARD_F_COMM_ERROR (_HRESULT_TYPEDEF_(0x80100013L))
value SCARD_F_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x80100001L))
value SCARD_F_UNKNOWN_ERROR (_HRESULT_TYPEDEF_(0x80100014L))
value SCARD_F_WAITED_TOO_LONG (_HRESULT_TYPEDEF_(0x80100007L))
value SCARD_LEAVE_CARD (0)
value SCARD_NEGOTIABLE (5)
value SCARD_POWERED (4)
value SCARD_POWER_DOWN (0)
value SCARD_PRESENT (2)
value SCARD_PROTOCOL_DEFAULT (0x80000000)
value SCARD_PROTOCOL_OPTIMAL (0x00000000)
value SCARD_PROTOCOL_RAW (0x00010000)
value SCARD_PROTOCOL_UNDEFINED (0x00000000)
value SCARD_PROVIDER_CSP (2)
value SCARD_PROVIDER_KSP (3)
value SCARD_PROVIDER_PRIMARY (1)
value SCARD_P_SHUTDOWN (_HRESULT_TYPEDEF_(0x80100018L))
value SCARD_READERSTATE_A (SCARD_READERSTATEA)
value SCARD_READERSTATE_W (SCARD_READERSTATEW)
value SCARD_READER_CONFISCATES (0x00000004)
value SCARD_READER_CONTACTLESS (0x00000008)
value SCARD_READER_EJECTS (0x00000002)
value SCARD_READER_SEL_AUTH_PACKAGE (((DWORD)-629))
value SCARD_READER_SWALLOWS (0x00000001)
value SCARD_READER_TYPE_EMBEDDEDSE (0x800)
value SCARD_READER_TYPE_IDE (0x10)
value SCARD_READER_TYPE_KEYBOARD (0x04)
value SCARD_READER_TYPE_NFC (0x100)
value SCARD_READER_TYPE_NGC (0x400)
value SCARD_READER_TYPE_PARALELL (0x02)
value SCARD_READER_TYPE_PCMCIA (0x40)
value SCARD_READER_TYPE_SCSI (0x08)
value SCARD_READER_TYPE_SERIAL (0x01)
value SCARD_READER_TYPE_TPM (0x80)
value SCARD_READER_TYPE_UICC (0x200)
value SCARD_READER_TYPE_USB (0x20)
value SCARD_READER_TYPE_VENDOR (0xF0)
value SCARD_RESET_CARD (1)
value SCARD_SCOPE_SYSTEM (2)
value SCARD_SCOPE_TERMINAL (1)
value SCARD_SCOPE_USER (0)
value SCARD_SHARE_DIRECT (3)
value SCARD_SHARE_EXCLUSIVE (1)
value SCARD_SHARE_SHARED (2)
value SCARD_SPECIFIC (6)
value SCARD_STATE_ATRMATCH (0x00000040)
value SCARD_STATE_CHANGED (0x00000002)
value SCARD_STATE_EMPTY (0x00000010)
value SCARD_STATE_EXCLUSIVE (0x00000080)
value SCARD_STATE_IGNORE (0x00000001)
value SCARD_STATE_INUSE (0x00000100)
value SCARD_STATE_MUTE (0x00000200)
value SCARD_STATE_PRESENT (0x00000020)
value SCARD_STATE_UNAVAILABLE (0x00000008)
value SCARD_STATE_UNAWARE (0x00000000)
value SCARD_STATE_UNKNOWN (0x00000004)
value SCARD_STATE_UNPOWERED (0x00000400)
value SCARD_SWALLOWED (3)
value SCARD_S_SUCCESS (NO_ERROR)
value SCARD_UNKNOWN (0)
value SCARD_UNPOWER_CARD (2)
value SCARD_WARM_RESET (2)
value SCARD_W_CACHE_ITEM_NOT_FOUND (_HRESULT_TYPEDEF_(0x80100070L))
value SCARD_W_CACHE_ITEM_STALE (_HRESULT_TYPEDEF_(0x80100071L))
value SCARD_W_CACHE_ITEM_TOO_BIG (_HRESULT_TYPEDEF_(0x80100072L))
value SCARD_W_CANCELLED_BY_USER (_HRESULT_TYPEDEF_(0x8010006EL))
value SCARD_W_CARD_NOT_AUTHENTICATED (_HRESULT_TYPEDEF_(0x8010006FL))
value SCARD_W_CHV_BLOCKED (_HRESULT_TYPEDEF_(0x8010006CL))
value SCARD_W_EOF (_HRESULT_TYPEDEF_(0x8010006DL))
value SCARD_W_REMOVED_CARD (_HRESULT_TYPEDEF_(0x80100069L))
value SCARD_W_RESET_CARD (_HRESULT_TYPEDEF_(0x80100068L))
value SCARD_W_SECURITY_VIOLATION (_HRESULT_TYPEDEF_(0x8010006AL))
value SCARD_W_UNPOWERED_CARD (_HRESULT_TYPEDEF_(0x80100067L))
value SCARD_W_UNRESPONSIVE_CARD (_HRESULT_TYPEDEF_(0x80100066L))
value SCARD_W_UNSUPPORTED_CARD (_HRESULT_TYPEDEF_(0x80100065L))
value SCARD_W_WRONG_CHV (_HRESULT_TYPEDEF_(0x8010006BL))
value SCERR_NOCARDNAME (0x4000)
value SCERR_NOGUIDS (0x8000)
value SCF_ISSECURE (0x00000001)
value SCHANNEL_ENC_KEY (0x00000001)
value SCHANNEL_MAC_KEY (0x00000000)
value SCHAR_MAX (127)
value SCHAR_MIN ((-128))
value SCHED_E_ACCOUNT_DBASE_CORRUPT (_HRESULT_TYPEDEF_(0x80041311L))
value SCHED_E_ACCOUNT_INFORMATION_NOT_SET (_HRESULT_TYPEDEF_(0x8004130FL))
value SCHED_E_ACCOUNT_NAME_NOT_FOUND (_HRESULT_TYPEDEF_(0x80041310L))
value SCHED_E_ALREADY_RUNNING (_HRESULT_TYPEDEF_(0x8004131FL))
value SCHED_E_CANNOT_OPEN_TASK (_HRESULT_TYPEDEF_(0x8004130DL))
value SCHED_E_DEPRECATED_FEATURE_USED (_HRESULT_TYPEDEF_(0x80041330L))
value SCHED_E_INVALIDVALUE (_HRESULT_TYPEDEF_(0x80041318L))
value SCHED_E_INVALID_TASK (_HRESULT_TYPEDEF_(0x8004130EL))
value SCHED_E_INVALID_TASK_HASH (_HRESULT_TYPEDEF_(0x80041321L))
value SCHED_E_MALFORMEDXML (_HRESULT_TYPEDEF_(0x8004131AL))
value SCHED_E_MISSINGNODE (_HRESULT_TYPEDEF_(0x80041319L))
value SCHED_E_NAMESPACE (_HRESULT_TYPEDEF_(0x80041317L))
value SCHED_E_NO_SECURITY_SERVICES (_HRESULT_TYPEDEF_(0x80041312L))
value SCHED_E_PAST_END_BOUNDARY (_HRESULT_TYPEDEF_(0x8004131EL))
value SCHED_E_SERVICE_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x80041322L))
value SCHED_E_SERVICE_NOT_INSTALLED (_HRESULT_TYPEDEF_(0x8004130CL))
value SCHED_E_SERVICE_NOT_LOCALSYSTEM (6200)
value SCHED_E_SERVICE_NOT_RUNNING (_HRESULT_TYPEDEF_(0x80041315L))
value SCHED_E_SERVICE_TOO_BUSY (_HRESULT_TYPEDEF_(0x80041323L))
value SCHED_E_START_ON_DEMAND (_HRESULT_TYPEDEF_(0x80041328L))
value SCHED_E_TASK_ATTEMPTED (_HRESULT_TYPEDEF_(0x80041324L))
value SCHED_E_TASK_DISABLED (_HRESULT_TYPEDEF_(0x80041326L))
value SCHED_E_TASK_NOT_READY (_HRESULT_TYPEDEF_(0x8004130AL))
value SCHED_E_TASK_NOT_RUNNING (_HRESULT_TYPEDEF_(0x8004130BL))
value SCHED_E_TASK_NOT_UBPM_COMPAT (_HRESULT_TYPEDEF_(0x80041329L))
value SCHED_E_TOO_MANY_NODES (_HRESULT_TYPEDEF_(0x8004131DL))
value SCHED_E_TRIGGER_NOT_FOUND (_HRESULT_TYPEDEF_(0x80041309L))
value SCHED_E_UNEXPECTEDNODE (_HRESULT_TYPEDEF_(0x80041316L))
value SCHED_E_UNKNOWN_OBJECT_VERSION (_HRESULT_TYPEDEF_(0x80041313L))
value SCHED_E_UNSUPPORTED_ACCOUNT_OPTION (_HRESULT_TYPEDEF_(0x80041314L))
value SCHED_E_USER_NOT_LOGGED_ON (_HRESULT_TYPEDEF_(0x80041320L))
value SCHED_S_BATCH_LOGON_PROBLEM (_HRESULT_TYPEDEF_(0x0004131CL))
value SCHED_S_EVENT_TRIGGER (_HRESULT_TYPEDEF_(0x00041308L))
value SCHED_S_SOME_TRIGGERS_FAILED (_HRESULT_TYPEDEF_(0x0004131BL))
value SCHED_S_TASK_DISABLED (_HRESULT_TYPEDEF_(0x00041302L))
value SCHED_S_TASK_HAS_NOT_RUN (_HRESULT_TYPEDEF_(0x00041303L))
value SCHED_S_TASK_NOT_SCHEDULED (_HRESULT_TYPEDEF_(0x00041305L))
value SCHED_S_TASK_NO_MORE_RUNS (_HRESULT_TYPEDEF_(0x00041304L))
value SCHED_S_TASK_NO_VALID_TRIGGERS (_HRESULT_TYPEDEF_(0x00041307L))
value SCHED_S_TASK_QUEUED (_HRESULT_TYPEDEF_(0x00041325L))
value SCHED_S_TASK_READY (_HRESULT_TYPEDEF_(0x00041300L))
value SCHED_S_TASK_RUNNING (_HRESULT_TYPEDEF_(0x00041301L))
value SCHED_S_TASK_TERMINATED (_HRESULT_TYPEDEF_(0x00041306L))
value SCM_MAX_SYMLINK_LEN_IN_CHARS (256)
value SCM_PD_FIRMWARE_LAST_DOWNLOAD (0x1)
value SCM_PD_FIRMWARE_REVISION_LENGTH_BYTES (32)
value SCM_PD_MAX_OPERATIONAL_STATUS (16)
value SCM_PD_MEMORY_SIZE_UNKNOWN (MAXDWORD64)
value SCM_PD_PROPERTY_NAME_LENGTH_IN_CHARS (128)
value SCM_REGION_SPA_UNKNOWN (MAXDWORD64)
value SCOPE_SECURITY_INFORMATION ((0x00000040L))
value SCREEN_FONTTYPE (0x2000)
value SCROLLLOCK_ON (0x0040)
value SCRUB_DATA_INPUT_FLAG_IGNORE_REDUNDANCY (0x00000008)
value SCRUB_DATA_INPUT_FLAG_OPLOCK_NOT_ACQUIRED (0x00000040)
value SCRUB_DATA_INPUT_FLAG_RESUME (0x00000001)
value SCRUB_DATA_INPUT_FLAG_SCRUB_BY_OBJECT_ID (0x00000020)
value SCRUB_DATA_INPUT_FLAG_SKIP_DATA (0x00000010)
value SCRUB_DATA_INPUT_FLAG_SKIP_IN_SYNC (0x00000002)
value SCRUB_DATA_INPUT_FLAG_SKIP_NON_INTEGRITY_DATA (0x00000004)
value SCRUB_DATA_OUTPUT_FLAG_INCOMPLETE (0x00000001)
value SCRUB_DATA_OUTPUT_FLAG_NON_USER_DATA_RANGE (0x00010000)
value SCRUB_DATA_OUTPUT_FLAG_PARITY_EXTENT_DATA_RETURNED (0x00020000)
value SCRUB_DATA_OUTPUT_FLAG_RESUME_CONTEXT_LENGTH_SPECIFIED (0x00040000)
value SCS_CAP_COMPSTR (0x00000001)
value SCS_CAP_MAKEREAD (0x00000002)
value SCS_CAP_SETRECONVERTSTRING (0x00000004)
value SCS_CHANGEATTR ((GCS_COMPREADATTR|GCS_COMPATTR))
value SCS_CHANGECLAUSE ((GCS_COMPREADCLAUSE|GCS_COMPCLAUSE))
value SCS_DOS_BINARY (1)
value SCS_PIF_BINARY (3)
value SCS_POSIX_BINARY (4)
value SCS_QUERYRECONVERTSTRING (0x00020000)
value SCS_SETRECONVERTSTRING (0x00010000)
value SCS_SETSTR ((GCS_COMPREADSTR|GCS_COMPSTR))
value SCS_THIS_PLATFORM_BINARY (SCS_64BIT_BINARY)
value SCS_WOW_BINARY (2)
value SC_ARRANGE (0xF110)
value SC_CLOSE (0xF060)
value SC_CONTEXTHELP (0xF180)
value SC_DEFAULT (0xF160)
value SC_DLG_FORCE_UI (0x04)
value SC_DLG_MINIMAL_UI (0x01)
value SC_DLG_NO_UI (0x02)
value SC_GROUP_IDENTIFIER (SC_GROUP_IDENTIFIERA)
value SC_HOTKEY (0xF150)
value SC_HSCROLL (0xF080)
value SC_ICON (SC_MINIMIZE)
value SC_KEYMENU (0xF100)
value SC_MANAGER_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | SC_MANAGER_CONNECT | SC_MANAGER_CREATE_SERVICE | SC_MANAGER_ENUMERATE_SERVICE | SC_MANAGER_LOCK | SC_MANAGER_QUERY_LOCK_STATUS | SC_MANAGER_MODIFY_BOOT_CONFIG))
value SC_MANAGER_CONNECT (0x0001)
value SC_MANAGER_CREATE_SERVICE (0x0002)
value SC_MANAGER_ENUMERATE_SERVICE (0x0004)
value SC_MANAGER_LOCK (0x0008)
value SC_MANAGER_MODIFY_BOOT_CONFIG (0x0020)
value SC_MANAGER_QUERY_LOCK_STATUS (0x0010)
value SC_MAXIMIZE (0xF030)
value SC_MINIMIZE (0xF020)
value SC_MONITORPOWER (0xF170)
value SC_MOUSEMENU (0xF090)
value SC_MOVE (0xF010)
value SC_NEXTWINDOW (0xF040)
value SC_PREVWINDOW (0xF050)
value SC_RESTORE (0xF120)
value SC_SCREENSAVE (0xF140)
value SC_SEPARATOR (0xF00F)
value SC_SIZE (0xF000)
value SC_TASKLIST (0xF130)
value SC_VSCROLL (0xF070)
value SC_ZOOM (SC_MAXIMIZE)
value SDC_ALLOW_CHANGES (0x00000400)
value SDC_ALLOW_PATH_ORDER_CHANGES (0x00002000)
value SDC_APPLY (0x00000080)
value SDC_FORCE_MODE_ENUMERATION (0x00001000)
value SDC_NO_OPTIMIZATION (0x00000100)
value SDC_PATH_PERSIST_IF_REQUIRED (0x00000800)
value SDC_SAVE_TO_DATABASE (0x00000200)
value SDC_TOPOLOGY_CLONE (0x00000002)
value SDC_TOPOLOGY_EXTEND (0x00000004)
value SDC_TOPOLOGY_EXTERNAL (0x00000008)
value SDC_TOPOLOGY_INTERNAL (0x00000001)
value SDC_TOPOLOGY_SUPPLIED (0x00000010)
value SDC_USE_DATABASE_CURRENT ((SDC_TOPOLOGY_INTERNAL | SDC_TOPOLOGY_CLONE | SDC_TOPOLOGY_EXTEND | SDC_TOPOLOGY_EXTERNAL))
value SDC_USE_SUPPLIED_DISPLAY_CONFIG (0x00000020)
value SDC_VALIDATE (0x00000040)
value SDC_VIRTUAL_MODE_AWARE (0x00008000)
value SDC_VIRTUAL_REFRESH_RATE_AWARE (0x00020000)
value SDIAG_E_CANCELLED (_NDIS_ERROR_TYPEDEF_(0x803C0100L))
value SDIAG_E_CANNOTRUN (_NDIS_ERROR_TYPEDEF_(0x803C0108L))
value SDIAG_E_DISABLED (_NDIS_ERROR_TYPEDEF_(0x803C0106L))
value SDIAG_E_MANAGEDHOST (_NDIS_ERROR_TYPEDEF_(0x803C0103L))
value SDIAG_E_NOVERIFIER (_NDIS_ERROR_TYPEDEF_(0x803C0104L))
value SDIAG_E_POWERSHELL (_NDIS_ERROR_TYPEDEF_(0x803C0102L))
value SDIAG_E_RESOURCE (_NDIS_ERROR_TYPEDEF_(0x803C010AL))
value SDIAG_E_ROOTCAUSE (_NDIS_ERROR_TYPEDEF_(0x803C010BL))
value SDIAG_E_SCRIPT (_NDIS_ERROR_TYPEDEF_(0x803C0101L))
value SDIAG_E_TRUST (_NDIS_ERROR_TYPEDEF_(0x803C0107L))
value SDIAG_E_VERSION (_NDIS_ERROR_TYPEDEF_(0x803C0109L))
value SDIAG_S_CANNOTRUN (_NDIS_ERROR_TYPEDEF_(0x003C0105L))
value SD_BOTH (0x02)
value SD_GLOBAL_CHANGE_TYPE_MACHINE_SID (1)
value SD_RECEIVE (0x00)
value SD_SEND (0x01)
value SEARCH_ALL (0x0)
value SEARCH_ALL_NO_SEQ (0x4)
value SEARCH_ALTERNATE (0x2)
value SEARCH_ALT_NO_SEQ (0x6)
value SEARCH_PRIMARY (0x1)
value SEARCH_PRI_NO_SEQ (0x5)
value SECTION_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED|SECTION_QUERY| SECTION_MAP_WRITE | SECTION_MAP_READ | SECTION_MAP_EXECUTE | SECTION_EXTEND_SIZE))
value SECTION_EXTEND_SIZE (0x0010)
value SECTION_MAP_EXECUTE (0x0008)
value SECTION_MAP_EXECUTE_EXPLICIT (0x0020)
value SECTION_MAP_READ (0x0004)
value SECTION_MAP_WRITE (0x0002)
value SECTION_QUERY (0x0001)
value SECURITY_ANONYMOUS_LOGON_RID ((0x00000007L))
value SECURITY_APPPOOL_ID_BASE_RID ((0x00000052L))
value SECURITY_APPPOOL_ID_RID_COUNT ((6L))
value SECURITY_APP_PACKAGE_BASE_RID ((0x00000002L))
value SECURITY_APP_PACKAGE_RID_COUNT ((8L))
value SECURITY_AUTHENTICATED_USER_RID ((0x0000000BL))
value SECURITY_AUTHENTICATION_AUTHORITY_ASSERTED_RID ((0x00000001L))
value SECURITY_AUTHENTICATION_AUTHORITY_RID_COUNT ((1L))
value SECURITY_AUTHENTICATION_FRESH_KEY_AUTH_RID ((0x00000003L))
value SECURITY_AUTHENTICATION_KEY_PROPERTY_ATTESTATION_RID ((0x00000006L))
value SECURITY_AUTHENTICATION_KEY_PROPERTY_MFA_RID ((0x00000005L))
value SECURITY_AUTHENTICATION_KEY_TRUST_RID ((0x00000004L))
value SECURITY_AUTHENTICATION_SERVICE_ASSERTED_RID ((0x00000002L))
value SECURITY_BATCH_RID ((0x00000003L))
value SECURITY_BUILTIN_APP_PACKAGE_RID_COUNT ((2L))
value SECURITY_BUILTIN_CAPABILITY_RID_COUNT ((2L))
value SECURITY_BUILTIN_DOMAIN_RID ((0x00000020L))
value SECURITY_BUILTIN_PACKAGE_ANY_PACKAGE ((0x00000001L))
value SECURITY_BUILTIN_PACKAGE_ANY_RESTRICTED_PACKAGE ((0x00000002L))
value SECURITY_CAPABILITY_APPOINTMENTS ((0x0000000BL))
value SECURITY_CAPABILITY_APP_RID ((0x00000400L))
value SECURITY_CAPABILITY_APP_SILO_RID ((0x00010000L))
value SECURITY_CAPABILITY_BASE_RID ((0x00000003L))
value SECURITY_CAPABILITY_CONTACTS ((0x0000000CL))
value SECURITY_CAPABILITY_DOCUMENTS_LIBRARY ((0x00000007L))
value SECURITY_CAPABILITY_ENTERPRISE_AUTHENTICATION ((0x00000008L))
value SECURITY_CAPABILITY_INTERNET_CLIENT ((0x00000001L))
value SECURITY_CAPABILITY_INTERNET_CLIENT_SERVER ((0x00000002L))
value SECURITY_CAPABILITY_INTERNET_EXPLORER ((0x00001000L))
value SECURITY_CAPABILITY_MUSIC_LIBRARY ((0x00000006L))
value SECURITY_CAPABILITY_PICTURES_LIBRARY ((0x00000004L))
value SECURITY_CAPABILITY_PRIVATE_NETWORK_CLIENT_SERVER ((0x00000003L))
value SECURITY_CAPABILITY_REMOVABLE_STORAGE ((0x0000000AL))
value SECURITY_CAPABILITY_RID_COUNT ((5L))
value SECURITY_CAPABILITY_SHARED_USER_CERTIFICATES ((0x00000009L))
value SECURITY_CAPABILITY_VIDEOS_LIBRARY ((0x00000005L))
value SECURITY_CCG_ID_BASE_RID ((0x0000005FL))
value SECURITY_CHILD_PACKAGE_RID_COUNT ((12L))
value SECURITY_CLOUD_INFRASTRUCTURE_SERVICES_ID_BASE_RID ((0x00000055L))
value SECURITY_CLOUD_INFRASTRUCTURE_SERVICES_ID_RID_COUNT ((6L))
value SECURITY_COM_ID_BASE_RID ((0x00000059L))
value SECURITY_CONTEXT_TRACKING (0x00040000)
value SECURITY_CREATOR_GROUP_RID ((0x00000001L))
value SECURITY_CREATOR_GROUP_SERVER_RID ((0x00000003L))
value SECURITY_CREATOR_OWNER_RID ((0x00000000L))
value SECURITY_CREATOR_OWNER_RIGHTS_RID ((0x00000004L))
value SECURITY_CREATOR_OWNER_SERVER_RID ((0x00000002L))
value SECURITY_CRED_TYPE_BASE_RID ((0x00000041L))
value SECURITY_CRED_TYPE_RID_COUNT ((2L))
value SECURITY_CRED_TYPE_THIS_ORG_CERT_RID ((0x00000001L))
value SECURITY_DASHOST_ID_BASE_RID ((0x0000005CL))
value SECURITY_DASHOST_ID_RID_COUNT ((6L))
value SECURITY_DESCRIPTOR_REVISION ((1))
value SECURITY_DIALUP_RID ((0x00000001L))
value SECURITY_DYNAMIC_TRACKING ((TRUE))
value SECURITY_EFFECTIVE_ONLY (0x00080000)
value SECURITY_ENTERPRISE_CONTROLLERS_RID ((0x00000009L))
value SECURITY_ENTERPRISE_READONLY_CONTROLLERS_RID ((0x00000016L))
value SECURITY_IE_STATE_GREEN (0x00000000)
value SECURITY_IE_STATE_RED (0x00000001)
value SECURITY_INSTALLER_CAPABILITY_RID_COUNT ((10))
value SECURITY_INSTALLER_GROUP_CAPABILITY_BASE ((0x20))
value SECURITY_INSTALLER_GROUP_CAPABILITY_RID_COUNT ((9))
value SECURITY_INTERACTIVE_RID ((0x00000004L))
value SECURITY_IUSER_RID ((0x00000011L))
value SECURITY_LOCAL_ACCOUNT_AND_ADMIN_RID ((0x00000072L))
value SECURITY_LOCAL_ACCOUNT_RID ((0x00000071L))
value SECURITY_LOCAL_LOGON_RID ((0x00000001L))
value SECURITY_LOCAL_RID ((0x00000000L))
value SECURITY_LOCAL_SERVICE_RID ((0x00000013L))
value SECURITY_LOCAL_SYSTEM_RID ((0x00000012L))
value SECURITY_LOGON_IDS_RID ((0x00000005L))
value SECURITY_LOGON_IDS_RID_COUNT ((3L))
value SECURITY_MANDATORY_HIGH_RID ((0x00003000L))
value SECURITY_MANDATORY_LOW_RID ((0x00001000L))
value SECURITY_MANDATORY_MAXIMUM_USER_RID (SECURITY_MANDATORY_SYSTEM_RID)
value SECURITY_MANDATORY_MEDIUM_PLUS_RID ((SECURITY_MANDATORY_MEDIUM_RID + 0x100))
value SECURITY_MANDATORY_MEDIUM_RID ((0x00002000L))
value SECURITY_MANDATORY_PROTECTED_PROCESS_RID ((0x00005000L))
value SECURITY_MANDATORY_SYSTEM_RID ((0x00004000L))
value SECURITY_MANDATORY_UNTRUSTED_RID ((0x00000000L))
value SECURITY_MAX_ALWAYS_FILTERED ((0x000003E7L))
value SECURITY_MAX_BASE_RID ((0x0000006FL))
value SECURITY_MIN_BASE_RID ((0x00000050L))
value SECURITY_MIN_NEVER_FILTERED ((0x000003E8L))
value SECURITY_NETWORK_RID ((0x00000002L))
value SECURITY_NETWORK_SERVICE_RID ((0x00000014L))
value SECURITY_NFS_ID_BASE_RID ((0x00000058L))
value SECURITY_NT_NON_UNIQUE ((0x00000015L))
value SECURITY_NT_NON_UNIQUE_SUB_AUTH_COUNT ((3L))
value SECURITY_NULL_RID ((0x00000000L))
value SECURITY_OTHER_ORGANIZATION_RID ((0x000003E8L))
value SECURITY_PACKAGE_BASE_RID ((0x00000040L))
value SECURITY_PACKAGE_DIGEST_RID ((0x00000015L))
value SECURITY_PACKAGE_NTLM_RID ((0x0000000AL))
value SECURITY_PACKAGE_RID_COUNT ((2L))
value SECURITY_PACKAGE_SCHANNEL_RID ((0x0000000EL))
value SECURITY_PARENT_PACKAGE_RID_COUNT ((SECURITY_APP_PACKAGE_RID_COUNT))
value SECURITY_PRINCIPAL_SELF_RID ((0x0000000AL))
value SECURITY_PROCESS_PROTECTION_LEVEL_ANTIMALWARE_RID ((0x00000600L))
value SECURITY_PROCESS_PROTECTION_LEVEL_APP_RID ((0x00000800L))
value SECURITY_PROCESS_PROTECTION_LEVEL_AUTHENTICODE_RID ((0x00000400L))
value SECURITY_PROCESS_PROTECTION_LEVEL_NONE_RID ((0x00000000L))
value SECURITY_PROCESS_PROTECTION_LEVEL_WINDOWS_RID ((0x00001000L))
value SECURITY_PROCESS_PROTECTION_LEVEL_WINTCB_RID ((0x00002000L))
value SECURITY_PROCESS_PROTECTION_TYPE_FULL_RID ((0x00000400L))
value SECURITY_PROCESS_PROTECTION_TYPE_LITE_RID ((0x00000200L))
value SECURITY_PROCESS_PROTECTION_TYPE_NONE_RID ((0x00000000L))
value SECURITY_PROCESS_TRUST_AUTHORITY_RID_COUNT ((2L))
value SECURITY_PROTOCOL_NONE (0x0000)
value SECURITY_PROXY_RID ((0x00000008L))
value SECURITY_RDV_GFX_BASE_RID ((0x0000005BL))
value SECURITY_REMOTE_LOGON_RID ((0x0000000EL))
value SECURITY_RESERVED_ID_BASE_RID ((0x00000051L))
value SECURITY_RESTRICTED_CODE_RID ((0x0000000CL))
value SECURITY_SERVER_LOGON_RID (SECURITY_ENTERPRISE_CONTROLLERS_RID)
value SECURITY_SERVICE_ID_BASE_RID ((0x00000050L))
value SECURITY_SERVICE_ID_RID_COUNT ((6L))
value SECURITY_SERVICE_RID ((0x00000006L))
value SECURITY_SQOS_PRESENT (0x00100000)
value SECURITY_STATIC_TRACKING ((FALSE))
value SECURITY_TASK_ID_BASE_RID ((0x00000057L))
value SECURITY_TERMINAL_SERVER_RID ((0x0000000DL))
value SECURITY_THIS_ORGANIZATION_RID ((0x0000000FL))
value SECURITY_UMFD_BASE_RID ((0x00000060L))
value SECURITY_USERMANAGER_ID_BASE_RID ((0x0000005DL))
value SECURITY_USERMANAGER_ID_RID_COUNT ((6L))
value SECURITY_USERMODEDRIVERHOST_ID_BASE_RID ((0x00000054L))
value SECURITY_USERMODEDRIVERHOST_ID_RID_COUNT ((6L))
value SECURITY_VALID_SQOS_FLAGS (0x001F0000)
value SECURITY_VIRTUALACCOUNT_ID_RID_COUNT ((6L))
value SECURITY_VIRTUALSERVER_ID_BASE_RID ((0x00000053L))
value SECURITY_VIRTUALSERVER_ID_RID_COUNT ((6L))
value SECURITY_WINDOWSMOBILE_ID_BASE_RID ((0x00000070L))
value SECURITY_WINDOW_MANAGER_BASE_RID ((0x0000005AL))
value SECURITY_WINRM_ID_BASE_RID ((0x0000005EL))
value SECURITY_WINRM_ID_RID_COUNT ((6L))
value SECURITY_WMIHOST_ID_BASE_RID ((0x00000056L))
value SECURITY_WMIHOST_ID_RID_COUNT ((6L))
value SECURITY_WORLD_RID ((0x00000000L))
value SECURITY_WRITE_RESTRICTED_CODE_RID ((0x00000021L))
value SEC_COMMIT (0x08000000)
value SEC_E_ALGORITHM_MISMATCH (_HRESULT_TYPEDEF_(0x80090331L))
value SEC_E_APPLICATION_PROTOCOL_MISMATCH (_HRESULT_TYPEDEF_(0x80090367L))
value SEC_E_BAD_BINDINGS (_HRESULT_TYPEDEF_(0x80090346L))
value SEC_E_BAD_PKGID (_HRESULT_TYPEDEF_(0x80090316L))
value SEC_E_BUFFER_TOO_SMALL (_HRESULT_TYPEDEF_(0x80090321L))
value SEC_E_CANNOT_INSTALL (_HRESULT_TYPEDEF_(0x80090307L))
value SEC_E_CANNOT_PACK (_HRESULT_TYPEDEF_(0x80090309L))
value SEC_E_CERT_EXPIRED (_HRESULT_TYPEDEF_(0x80090328L))
value SEC_E_CERT_UNKNOWN (_HRESULT_TYPEDEF_(0x80090327L))
value SEC_E_CERT_WRONG_USAGE (_HRESULT_TYPEDEF_(0x80090349L))
value SEC_E_CONTEXT_EXPIRED (_HRESULT_TYPEDEF_(0x80090317L))
value SEC_E_CROSSREALM_DELEGATION_FAILURE (_HRESULT_TYPEDEF_(0x80090357L))
value SEC_E_CRYPTO_SYSTEM_INVALID (_HRESULT_TYPEDEF_(0x80090337L))
value SEC_E_DECRYPT_FAILURE (_HRESULT_TYPEDEF_(0x80090330L))
value SEC_E_DELEGATION_POLICY (_HRESULT_TYPEDEF_(0x8009035EL))
value SEC_E_DELEGATION_REQUIRED (_HRESULT_TYPEDEF_(0x80090345L))
value SEC_E_DOWNGRADE_DETECTED (_HRESULT_TYPEDEF_(0x80090350L))
value SEC_E_ENCRYPT_FAILURE (_HRESULT_TYPEDEF_(0x80090329L))
value SEC_E_EXT_BUFFER_TOO_SMALL (_HRESULT_TYPEDEF_(0x8009036AL))
value SEC_E_ILLEGAL_MESSAGE (_HRESULT_TYPEDEF_(0x80090326L))
value SEC_E_INCOMPLETE_CREDENTIALS (_HRESULT_TYPEDEF_(0x80090320L))
value SEC_E_INCOMPLETE_MESSAGE (_HRESULT_TYPEDEF_(0x80090318L))
value SEC_E_INSUFFICIENT_BUFFERS (_HRESULT_TYPEDEF_(0x8009036BL))
value SEC_E_INSUFFICIENT_MEMORY (_HRESULT_TYPEDEF_(0x80090300L))
value SEC_E_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x80090304L))
value SEC_E_INVALID_HANDLE (_HRESULT_TYPEDEF_(0x80090301L))
value SEC_E_INVALID_PARAMETER (_HRESULT_TYPEDEF_(0x8009035DL))
value SEC_E_INVALID_TOKEN (_HRESULT_TYPEDEF_(0x80090308L))
value SEC_E_INVALID_UPN_NAME (_HRESULT_TYPEDEF_(0x80090369L))
value SEC_E_ISSUING_CA_UNTRUSTED (_HRESULT_TYPEDEF_(0x80090352L))
value SEC_E_ISSUING_CA_UNTRUSTED_KDC (_HRESULT_TYPEDEF_(0x80090359L))
value SEC_E_KDC_CERT_EXPIRED (_HRESULT_TYPEDEF_(0x8009035AL))
value SEC_E_KDC_CERT_REVOKED (_HRESULT_TYPEDEF_(0x8009035BL))
value SEC_E_KDC_INVALID_REQUEST (_HRESULT_TYPEDEF_(0x80090340L))
value SEC_E_KDC_UNABLE_TO_REFER (_HRESULT_TYPEDEF_(0x80090341L))
value SEC_E_KDC_UNKNOWN_ETYPE (_HRESULT_TYPEDEF_(0x80090342L))
value SEC_E_LOGON_DENIED (_HRESULT_TYPEDEF_(0x8009030CL))
value SEC_E_MAX_REFERRALS_EXCEEDED (_HRESULT_TYPEDEF_(0x80090338L))
value SEC_E_MESSAGE_ALTERED (_HRESULT_TYPEDEF_(0x8009030FL))
value SEC_E_MULTIPLE_ACCOUNTS (_HRESULT_TYPEDEF_(0x80090347L))
value SEC_E_MUST_BE_KDC (_HRESULT_TYPEDEF_(0x80090339L))
value SEC_E_MUTUAL_AUTH_FAILED (_HRESULT_TYPEDEF_(0x80090363L))
value SEC_E_NOT_OWNER (_HRESULT_TYPEDEF_(0x80090306L))
value SEC_E_NOT_SUPPORTED (SEC_E_UNSUPPORTED_FUNCTION)
value SEC_E_NO_AUTHENTICATING_AUTHORITY (_HRESULT_TYPEDEF_(0x80090311L))
value SEC_E_NO_CONTEXT (_HRESULT_TYPEDEF_(0x80090361L))
value SEC_E_NO_CREDENTIALS (_HRESULT_TYPEDEF_(0x8009030EL))
value SEC_E_NO_IMPERSONATION (_HRESULT_TYPEDEF_(0x8009030BL))
value SEC_E_NO_IP_ADDRESSES (_HRESULT_TYPEDEF_(0x80090335L))
value SEC_E_NO_KERB_KEY (_HRESULT_TYPEDEF_(0x80090348L))
value SEC_E_NO_PA_DATA (_HRESULT_TYPEDEF_(0x8009033CL))
value SEC_E_NO_SPM (SEC_E_INTERNAL_ERROR)
value SEC_E_NO_TGT_REPLY (_HRESULT_TYPEDEF_(0x80090334L))
value SEC_E_OK (((HRESULT)0x00000000L))
value SEC_E_ONLY_HTTPS_ALLOWED (_HRESULT_TYPEDEF_(0x80090365L))
value SEC_E_OUT_OF_SEQUENCE (_HRESULT_TYPEDEF_(0x80090310L))
value SEC_E_PKINIT_CLIENT_FAILURE (_HRESULT_TYPEDEF_(0x80090354L))
value SEC_E_PKINIT_NAME_MISMATCH (_HRESULT_TYPEDEF_(0x8009033DL))
value SEC_E_POLICY_NLTM_ONLY (_HRESULT_TYPEDEF_(0x8009035FL))
value SEC_E_QOP_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8009030AL))
value SEC_E_REVOCATION_OFFLINE_C (_HRESULT_TYPEDEF_(0x80090353L))
value SEC_E_REVOCATION_OFFLINE_KDC (_HRESULT_TYPEDEF_(0x80090358L))
value SEC_E_SECPKG_NOT_FOUND (_HRESULT_TYPEDEF_(0x80090305L))
value SEC_E_SECURITY_QOS_FAILED (_HRESULT_TYPEDEF_(0x80090332L))
value SEC_E_SHUTDOWN_IN_PROGRESS (_HRESULT_TYPEDEF_(0x8009033FL))
value SEC_E_SMARTCARD_CERT_EXPIRED (_HRESULT_TYPEDEF_(0x80090355L))
value SEC_E_SMARTCARD_CERT_REVOKED (_HRESULT_TYPEDEF_(0x80090351L))
value SEC_E_SMARTCARD_LOGON_REQUIRED (_HRESULT_TYPEDEF_(0x8009033EL))
value SEC_E_STRONG_CRYPTO_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8009033AL))
value SEC_E_TARGET_UNKNOWN (_HRESULT_TYPEDEF_(0x80090303L))
value SEC_E_TIME_SKEW (_HRESULT_TYPEDEF_(0x80090324L))
value SEC_E_TOO_MANY_PRINCIPALS (_HRESULT_TYPEDEF_(0x8009033BL))
value SEC_E_UNFINISHED_CONTEXT_DELETED (_HRESULT_TYPEDEF_(0x80090333L))
value SEC_E_UNKNOWN_CREDENTIALS (_HRESULT_TYPEDEF_(0x8009030DL))
value SEC_E_UNSUPPORTED_FUNCTION (_HRESULT_TYPEDEF_(0x80090302L))
value SEC_E_UNSUPPORTED_PREAUTH (_HRESULT_TYPEDEF_(0x80090343L))
value SEC_E_UNTRUSTED_ROOT (_HRESULT_TYPEDEF_(0x80090325L))
value SEC_E_WRONG_CREDENTIAL_HANDLE (_HRESULT_TYPEDEF_(0x80090336L))
value SEC_E_WRONG_PRINCIPAL (_HRESULT_TYPEDEF_(0x80090322L))
value SEC_FILE (0x00800000)
value SEC_HUGE_PAGES (0x00020000)
value SEC_IMAGE (0x01000000)
value SEC_IMAGE_NO_EXECUTE ((SEC_IMAGE | SEC_NOCACHE))
value SEC_I_ASYNC_CALL_PENDING (_HRESULT_TYPEDEF_(0x00090368L))
value SEC_I_COMPLETE_AND_CONTINUE (_HRESULT_TYPEDEF_(0x00090314L))
value SEC_I_COMPLETE_NEEDED (_HRESULT_TYPEDEF_(0x00090313L))
value SEC_I_CONTEXT_EXPIRED (_HRESULT_TYPEDEF_(0x00090317L))
value SEC_I_CONTINUE_NEEDED (_HRESULT_TYPEDEF_(0x00090312L))
value SEC_I_CONTINUE_NEEDED_MESSAGE_OK (_HRESULT_TYPEDEF_(0x00090366L))
value SEC_I_GENERIC_EXTENSION_RECEIVED (_HRESULT_TYPEDEF_(0x00090316L))
value SEC_I_INCOMPLETE_CREDENTIALS (_HRESULT_TYPEDEF_(0x00090320L))
value SEC_I_LOCAL_LOGON (_HRESULT_TYPEDEF_(0x00090315L))
value SEC_I_MESSAGE_FRAGMENT (_HRESULT_TYPEDEF_(0x00090364L))
value SEC_I_NO_LSA_CONTEXT (_HRESULT_TYPEDEF_(0x00090323L))
value SEC_I_NO_RENEGOTIATION (_HRESULT_TYPEDEF_(0x00090360L))
value SEC_I_RENEGOTIATE (_HRESULT_TYPEDEF_(0x00090321L))
value SEC_I_SIGNATURE_NEEDED (_HRESULT_TYPEDEF_(0x0009035CL))
value SEC_LARGE_PAGES (0x80000000)
value SEC_NOCACHE (0x10000000)
value SEC_PARTITION_OWNER_HANDLE (0x00040000)
value SEC_PROTECTED_IMAGE (0x02000000)
value SEC_RESERVE (0x04000000)
value SEC_WINNT_AUTH_IDENTITY (SEC_WINNT_AUTH_IDENTITY_A)
value SEC_WINNT_AUTH_IDENTITY_ANSI (0x1)
value SEC_WINNT_AUTH_IDENTITY_UNICODE (0x2)
value SEC_WRITECOMBINE (0x40000000)
value SEEK_CUR (1)
value SEEK_END (2)
value SEEK_SET (0)
value SEE_MASK_ASYNCOK (0x00100000)
value SEE_MASK_CLASSKEY (0x00000003)
value SEE_MASK_CLASSNAME (0x00000001)
value SEE_MASK_CONNECTNETDRV (0x00000080)
value SEE_MASK_DEFAULT (0x00000000)
value SEE_MASK_DOENVSUBST (0x00000200)
value SEE_MASK_FLAG_DDEWAIT (SEE_MASK_NOASYNC)
value SEE_MASK_FLAG_HINST_IS_SITE (0x08000000)
value SEE_MASK_FLAG_LOG_USAGE (0x04000000)
value SEE_MASK_FLAG_NO_UI (0x00000400)
value SEE_MASK_HMONITOR (0x00200000)
value SEE_MASK_HOTKEY (0x00000020)
value SEE_MASK_IDLIST (0x00000004)
value SEE_MASK_INVOKEIDLIST (0x0000000c)
value SEE_MASK_NOASYNC (0x00000100)
value SEE_MASK_NOCLOSEPROCESS (0x00000040)
value SEE_MASK_NOQUERYCLASSSTORE (0x01000000)
value SEE_MASK_NOZONECHECKS (0x00800000)
value SEE_MASK_NO_CONSOLE (0x00008000)
value SEE_MASK_UNICODE (0x00004000)
value SEE_MASK_WAITFORINPUTIDLE (0x02000000)
value SEF_AI_USE_EXTRA_PARAMS (0x800)
value SEF_AVOID_OWNER_CHECK (0x10)
value SEF_AVOID_OWNER_RESTRICTION (0x1000)
value SEF_AVOID_PRIVILEGE_CHECK (0x08)
value SEF_DACL_AUTO_INHERIT (0x01)
value SEF_DEFAULT_DESCRIPTOR_FOR_OBJECT (0x04)
value SEF_DEFAULT_GROUP_FROM_PARENT (0x40)
value SEF_DEFAULT_OWNER_FROM_PARENT (0x20)
value SEF_FORCE_USER_MODE (0x2000)
value SEF_MACL_NO_EXECUTE_UP (0x400)
value SEF_MACL_NO_READ_UP (0x200)
value SEF_MACL_NO_WRITE_UP (0x100)
value SEF_MACL_VALID_FLAGS ((SEF_MACL_NO_WRITE_UP | SEF_MACL_NO_READ_UP | SEF_MACL_NO_EXECUTE_UP))
value SEF_NORMALIZE_OUTPUT_DESCRIPTOR (0x4000)
value SEF_SACL_AUTO_INHERIT (0x02)
value SELECTDIB (41)
value SELECTPAPERSOURCE (18)
value SELECT_CAP_CONVERSION (0x00000001)
value SELECT_CAP_SENTENCE (0x00000002)
value SEMAPHORE_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED|SYNCHRONIZE|0x3))
value SEMAPHORE_MODIFY_STATE (0x0002)
value SEM_FAILCRITICALERRORS (0x0001)
value SEM_NOALIGNMENTFAULTEXCEPT (0x0004)
value SEM_NOGPFAULTERRORBOX (0x0002)
value SEM_NOOPENFILEERRORBOX (0x8000)
value SERIAL_IOC_FCR_DMA_MODE (((DWORD)0x00000008))
value SERIAL_IOC_FCR_FIFO_ENABLE (((DWORD)0x00000001))
value SERIAL_IOC_FCR_RCVR_RESET (((DWORD)0x00000002))
value SERIAL_IOC_FCR_RCVR_TRIGGER_LSB (((DWORD)0x00000040))
value SERIAL_IOC_FCR_RCVR_TRIGGER_MSB (((DWORD)0x00000080))
value SERIAL_IOC_FCR_XMIT_RESET (((DWORD)0x00000004))
value SERIAL_IOC_MCR_DTR (((DWORD)0x00000001))
value SERIAL_IOC_MCR_LOOP (((DWORD)0x00000010))
value SERIAL_IOC_MCR_RTS (((DWORD)0x00000002))
value SERIAL_LSRMST_ESCAPE (((BYTE )0x00))
value SERIAL_LSRMST_LSR_DATA (((BYTE )0x01))
value SERIAL_LSRMST_LSR_NODATA (((BYTE )0x02))
value SERIAL_LSRMST_MST (((BYTE )0x03))
value SERIAL_NUMBER_LENGTH (32)
value SERKF_AVAILABLE (0x00000002)
value SERKF_INDICATOR (0x00000004)
value SERKF_SERIALKEYSON (0x00000001)
value SERVER_ACCESS_ADMINISTER (0x00000001)
value SERVER_ACCESS_ENUMERATE (0x00000002)
value SERVER_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | SERVER_ACCESS_ADMINISTER | SERVER_ACCESS_ENUMERATE))
value SERVER_EXECUTE ((STANDARD_RIGHTS_EXECUTE | SERVER_ACCESS_ENUMERATE))
value SERVER_NOTIFY_FIELD_PRINT_DRIVER_ISOLATION_GROUP (0x00)
value SERVER_NOTIFY_TYPE (0x02)
value SERVER_READ ((STANDARD_RIGHTS_READ | SERVER_ACCESS_ENUMERATE))
value SERVER_WRITE ((STANDARD_RIGHTS_WRITE | SERVER_ACCESS_ADMINISTER | SERVER_ACCESS_ENUMERATE))
value SERVICES_ACTIVE_DATABASE (SERVICES_ACTIVE_DATABASEA)
value SERVICES_FAILED_DATABASE (SERVICES_FAILED_DATABASEA)
value SERVICETYPE_BESTEFFORT (0x00000001)
value SERVICETYPE_CONTROLLEDLOAD (0x00000002)
value SERVICETYPE_GENERAL_INFORMATION (0x00000005)
value SERVICETYPE_GUARANTEED (0x00000003)
value SERVICETYPE_NETWORK_CONTROL (0x0000000A)
value SERVICETYPE_NETWORK_UNAVAILABLE (0x00000004)
value SERVICETYPE_NOCHANGE (0x00000006)
value SERVICETYPE_NONCONFORMING (0x00000009)
value SERVICETYPE_NOTRAFFIC (0x00000000)
value SERVICETYPE_QUALITATIVE (0x0000000D)
value SERVICE_ACCEPT_HARDWAREPROFILECHANGE (0x00000020)
value SERVICE_ACCEPT_LOWRESOURCES (0x00002000)
value SERVICE_ACCEPT_NETBINDCHANGE (0x00000010)
value SERVICE_ACCEPT_PARAMCHANGE (0x00000008)
value SERVICE_ACCEPT_PAUSE_CONTINUE (0x00000002)
value SERVICE_ACCEPT_POWEREVENT (0x00000040)
value SERVICE_ACCEPT_PRESHUTDOWN (0x00000100)
value SERVICE_ACCEPT_SESSIONCHANGE (0x00000080)
value SERVICE_ACCEPT_SHUTDOWN (0x00000004)
value SERVICE_ACCEPT_STOP (0x00000001)
value SERVICE_ACCEPT_SYSTEMLOWRESOURCES (0x00004000)
value SERVICE_ACCEPT_TIMECHANGE (0x00000200)
value SERVICE_ACCEPT_TRIGGEREVENT (0x00000400)
value SERVICE_ACCEPT_USER_LOGOFF (0x00000800)
value SERVICE_ACTIVE (0x00000001)
value SERVICE_ADAPTER (0x00000004)
value SERVICE_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | SERVICE_QUERY_CONFIG | SERVICE_CHANGE_CONFIG | SERVICE_QUERY_STATUS | SERVICE_ENUMERATE_DEPENDENTS | SERVICE_START | SERVICE_STOP | SERVICE_PAUSE_CONTINUE | SERVICE_INTERROGATE | SERVICE_USER_DEFINED_CONTROL))
value SERVICE_AUTO_START (0x00000002)
value SERVICE_BESTEFFORT (0x80010000)
value SERVICE_BOOT_START (0x00000000)
value SERVICE_CHANGE_CONFIG (0x0002)
value SERVICE_CONFIG_DELAYED_AUTO_START_INFO (3)
value SERVICE_CONFIG_DESCRIPTION (1)
value SERVICE_CONFIG_FAILURE_ACTIONS (2)
value SERVICE_CONFIG_FAILURE_ACTIONS_FLAG (4)
value SERVICE_CONFIG_LAUNCH_PROTECTED (12)
value SERVICE_CONFIG_PREFERRED_NODE (9)
value SERVICE_CONFIG_PRESHUTDOWN_INFO (7)
value SERVICE_CONFIG_REQUIRED_PRIVILEGES_INFO (6)
value SERVICE_CONFIG_SERVICE_SID_INFO (5)
value SERVICE_CONFIG_TRIGGER_INFO (8)
value SERVICE_CONTINUE_PENDING (0x00000005)
value SERVICE_CONTROLLEDLOAD (0x80020000)
value SERVICE_CONTROL_CONTINUE (0x00000003)
value SERVICE_CONTROL_DEVICEEVENT (0x0000000B)
value SERVICE_CONTROL_HARDWAREPROFILECHANGE (0x0000000C)
value SERVICE_CONTROL_INTERROGATE (0x00000004)
value SERVICE_CONTROL_LOWRESOURCES (0x00000060)
value SERVICE_CONTROL_NETBINDADD (0x00000007)
value SERVICE_CONTROL_NETBINDDISABLE (0x0000000A)
value SERVICE_CONTROL_NETBINDENABLE (0x00000009)
value SERVICE_CONTROL_NETBINDREMOVE (0x00000008)
value SERVICE_CONTROL_PARAMCHANGE (0x00000006)
value SERVICE_CONTROL_PAUSE (0x00000002)
value SERVICE_CONTROL_POWEREVENT (0x0000000D)
value SERVICE_CONTROL_PRESHUTDOWN (0x0000000F)
value SERVICE_CONTROL_SESSIONCHANGE (0x0000000E)
value SERVICE_CONTROL_SHUTDOWN (0x00000005)
value SERVICE_CONTROL_STATUS_REASON_INFO (1)
value SERVICE_CONTROL_STOP (0x00000001)
value SERVICE_CONTROL_SYSTEMLOWRESOURCES (0x00000061)
value SERVICE_CONTROL_TIMECHANGE (0x00000010)
value SERVICE_CONTROL_TRIGGEREVENT (0x00000020)
value SERVICE_DEMAND_START (0x00000003)
value SERVICE_DISABLED (0x00000004)
value SERVICE_DRIVER ((SERVICE_KERNEL_DRIVER | SERVICE_FILE_SYSTEM_DRIVER | SERVICE_RECOGNIZER_DRIVER))
value SERVICE_DYNAMIC_INFORMATION_LEVEL_START_REASON (1)
value SERVICE_ENUMERATE_DEPENDENTS (0x0008)
value SERVICE_ERROR_CRITICAL (0x00000003)
value SERVICE_ERROR_IGNORE (0x00000000)
value SERVICE_ERROR_NORMAL (0x00000001)
value SERVICE_ERROR_SEVERE (0x00000002)
value SERVICE_FILE_SYSTEM_DRIVER (0x00000002)
value SERVICE_GUARANTEED (0x80040000)
value SERVICE_INACTIVE (0x00000002)
value SERVICE_INTERACTIVE_PROCESS (0x00000100)
value SERVICE_INTERROGATE (0x0080)
value SERVICE_KERNEL_DRIVER (0x00000001)
value SERVICE_LAUNCH_PROTECTED_ANTIMALWARE_LIGHT (3)
value SERVICE_LAUNCH_PROTECTED_NONE (0)
value SERVICE_LAUNCH_PROTECTED_WINDOWS (1)
value SERVICE_LAUNCH_PROTECTED_WINDOWS_LIGHT (2)
value SERVICE_MAIN_FUNCTION (SERVICE_MAIN_FUNCTIONA)
value SERVICE_MULTIPLE ((0x00000001))
value SERVICE_NOTIFY_CONTINUE_PENDING (0x00000010)
value SERVICE_NOTIFY_CREATED (0x00000080)
value SERVICE_NOTIFY_DELETED (0x00000100)
value SERVICE_NOTIFY_DELETE_PENDING (0x00000200)
value SERVICE_NOTIFY_PAUSED (0x00000040)
value SERVICE_NOTIFY_PAUSE_PENDING (0x00000020)
value SERVICE_NOTIFY_RUNNING (0x00000008)
value SERVICE_NOTIFY_START_PENDING (0x00000002)
value SERVICE_NOTIFY_STATUS_CHANGE (SERVICE_NOTIFY_STATUS_CHANGE_2)
value SERVICE_NOTIFY_STOPPED (0x00000001)
value SERVICE_NOTIFY_STOP_PENDING (0x00000004)
value SERVICE_NO_CHANGE (0xffffffff)
value SERVICE_NO_QOS_SIGNALING (0x40000000)
value SERVICE_NO_TRAFFIC_CONTROL (0x81000000)
value SERVICE_PAUSED (0x00000007)
value SERVICE_PAUSE_CONTINUE (0x0040)
value SERVICE_PAUSE_PENDING (0x00000006)
value SERVICE_PKG_SERVICE (0x00000200)
value SERVICE_QUALITATIVE (0x80200000)
value SERVICE_QUERY_CONFIG (0x0001)
value SERVICE_QUERY_STATUS (0x0004)
value SERVICE_RECOGNIZER_DRIVER (0x00000008)
value SERVICE_RUNNING (0x00000004)
value SERVICE_RUNS_IN_SYSTEM_PROCESS (0x00000001)
value SERVICE_SID_TYPE_NONE (0x00000000)
value SERVICE_SID_TYPE_RESTRICTED (( 0x00000002 | SERVICE_SID_TYPE_UNRESTRICTED ))
value SERVICE_SID_TYPE_UNRESTRICTED (0x00000001)
value SERVICE_START (0x0010)
value SERVICE_START_PENDING (0x00000002)
value SERVICE_START_REASON_AUTO (0x00000002)
value SERVICE_START_REASON_DELAYEDAUTO (0x00000010)
value SERVICE_START_REASON_DEMAND (0x00000001)
value SERVICE_START_REASON_RESTART_ON_FAILURE (0x00000008)
value SERVICE_START_REASON_TRIGGER (0x00000004)
value SERVICE_STATE_ALL ((SERVICE_ACTIVE | SERVICE_INACTIVE))
value SERVICE_STOP (0x0020)
value SERVICE_STOPPED (0x00000001)
value SERVICE_STOP_PENDING (0x00000003)
value SERVICE_STOP_REASON_FLAG_CUSTOM (0x20000000)
value SERVICE_STOP_REASON_FLAG_MAX (0x80000000)
value SERVICE_STOP_REASON_FLAG_MIN (0x00000000)
value SERVICE_STOP_REASON_FLAG_PLANNED (0x40000000)
value SERVICE_STOP_REASON_FLAG_UNPLANNED (0x10000000)
value SERVICE_STOP_REASON_MAJOR_APPLICATION (0x00050000)
value SERVICE_STOP_REASON_MAJOR_HARDWARE (0x00020000)
value SERVICE_STOP_REASON_MAJOR_MAX (0x00070000)
value SERVICE_STOP_REASON_MAJOR_MAX_CUSTOM (0x00ff0000)
value SERVICE_STOP_REASON_MAJOR_MIN (0x00000000)
value SERVICE_STOP_REASON_MAJOR_MIN_CUSTOM (0x00400000)
value SERVICE_STOP_REASON_MAJOR_NONE (0x00060000)
value SERVICE_STOP_REASON_MAJOR_OPERATINGSYSTEM (0x00030000)
value SERVICE_STOP_REASON_MAJOR_OTHER (0x00010000)
value SERVICE_STOP_REASON_MAJOR_SOFTWARE (0x00040000)
value SERVICE_STOP_REASON_MINOR_DISK (0x00000008)
value SERVICE_STOP_REASON_MINOR_ENVIRONMENT (0x0000000a)
value SERVICE_STOP_REASON_MINOR_HARDWARE_DRIVER (0x0000000b)
value SERVICE_STOP_REASON_MINOR_HUNG (0x00000006)
value SERVICE_STOP_REASON_MINOR_INSTALLATION (0x00000003)
value SERVICE_STOP_REASON_MINOR_MAINTENANCE (0x00000002)
value SERVICE_STOP_REASON_MINOR_MAX (0x00000019)
value SERVICE_STOP_REASON_MINOR_MAX_CUSTOM (0x0000FFFF)
value SERVICE_STOP_REASON_MINOR_MEMOTYLIMIT (0x00000018)
value SERVICE_STOP_REASON_MINOR_MIN (0x00000000)
value SERVICE_STOP_REASON_MINOR_MIN_CUSTOM (0x00000100)
value SERVICE_STOP_REASON_MINOR_MMC (0x00000016)
value SERVICE_STOP_REASON_MINOR_NETWORKCARD (0x00000009)
value SERVICE_STOP_REASON_MINOR_NETWORK_CONNECTIVITY (0x00000011)
value SERVICE_STOP_REASON_MINOR_NONE (0x00000017)
value SERVICE_STOP_REASON_MINOR_OTHER (0x00000001)
value SERVICE_STOP_REASON_MINOR_OTHERDRIVER (0x0000000c)
value SERVICE_STOP_REASON_MINOR_RECONFIG (0x00000005)
value SERVICE_STOP_REASON_MINOR_SECURITY (0x00000010)
value SERVICE_STOP_REASON_MINOR_SECURITYFIX (0x0000000f)
value SERVICE_STOP_REASON_MINOR_SECURITYFIX_UNINSTALL (0x00000015)
value SERVICE_STOP_REASON_MINOR_SERVICEPACK (0x0000000d)
value SERVICE_STOP_REASON_MINOR_SERVICEPACK_UNINSTALL (0x00000013)
value SERVICE_STOP_REASON_MINOR_SOFTWARE_UPDATE (0x0000000e)
value SERVICE_STOP_REASON_MINOR_SOFTWARE_UPDATE_UNINSTALL (0x00000014)
value SERVICE_STOP_REASON_MINOR_UNSTABLE (0x00000007)
value SERVICE_STOP_REASON_MINOR_UPGRADE (0x00000004)
value SERVICE_STOP_REASON_MINOR_WMI (0x00000012)
value SERVICE_SYSTEM_START (0x00000001)
value SERVICE_TRIGGER_ACTION_SERVICE_START (1)
value SERVICE_TRIGGER_ACTION_SERVICE_STOP (2)
value SERVICE_TRIGGER_DATA_TYPE_BINARY (1)
value SERVICE_TRIGGER_DATA_TYPE_KEYWORD_ALL (5)
value SERVICE_TRIGGER_DATA_TYPE_KEYWORD_ANY (4)
value SERVICE_TRIGGER_DATA_TYPE_LEVEL (3)
value SERVICE_TRIGGER_DATA_TYPE_STRING (2)
value SERVICE_TRIGGER_TYPE_AGGREGATE (30)
value SERVICE_TRIGGER_TYPE_CUSTOM (20)
value SERVICE_TRIGGER_TYPE_CUSTOM_SYSTEM_STATE_CHANGE (7)
value SERVICE_TRIGGER_TYPE_DEVICE_INTERFACE_ARRIVAL (1)
value SERVICE_TRIGGER_TYPE_DOMAIN_JOIN (3)
value SERVICE_TRIGGER_TYPE_FIREWALL_PORT_EVENT (4)
value SERVICE_TRIGGER_TYPE_GROUP_POLICY (5)
value SERVICE_TRIGGER_TYPE_IP_ADDRESS_AVAILABILITY (2)
value SERVICE_TRIGGER_TYPE_NETWORK_ENDPOINT (6)
value SERVICE_TYPE_ALL ((SERVICE_WIN32 | SERVICE_ADAPTER | SERVICE_DRIVER | SERVICE_INTERACTIVE_PROCESS | SERVICE_USER_SERVICE | SERVICE_USERSERVICE_INSTANCE | SERVICE_PKG_SERVICE))
value SERVICE_TYPE_VALUE_OBJECTID (SERVICE_TYPE_VALUE_OBJECTIDA)
value SERVICE_TYPE_VALUE_SAPID (SERVICE_TYPE_VALUE_SAPIDA)
value SERVICE_TYPE_VALUE_TCPPORT (SERVICE_TYPE_VALUE_TCPPORTA)
value SERVICE_TYPE_VALUE_UDPPORT (SERVICE_TYPE_VALUE_UDPPORTA)
value SERVICE_USERSERVICE_INSTANCE (0x00000080)
value SERVICE_USER_DEFINED_CONTROL (0x0100)
value SERVICE_USER_OWN_PROCESS ((SERVICE_USER_SERVICE | SERVICE_WIN32_OWN_PROCESS))
value SERVICE_USER_SERVICE (0x00000040)
value SERVICE_USER_SHARE_PROCESS ((SERVICE_USER_SERVICE | SERVICE_WIN32_SHARE_PROCESS))
value SESSION_ABORTED (0x06)
value SESSION_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | SESSION_QUERY_ACCESS | SESSION_MODIFY_ACCESS))
value SESSION_ESTABLISHED (0x03)
value SESSION_MODIFY_ACCESS (0x0002)
value SESSION_QUERY_ACCESS (0x0001)
value SETABORTPROC (9)
value SETALLJUSTVALUES (771)
value SETBREAK (8)
value SETCHARSET (772)
value SETCOLORTABLE (4)
value SETCOPYCOUNT (17)
value SETDIBSCALING (32)
value SETDTR (5)
value SETICMPROFILE_EMBEDED (0x00000001)
value SETKERNTRACK (770)
value SETLINECAP (21)
value SETLINEJOIN (22)
value SETMITERLIMIT (23)
value SETRGBSTRING (SETRGBSTRINGA)
value SETRTS (3)
value SETWALLPAPER_DEFAULT (((LPWSTR)-1))
value SETXOFF (1)
value SETXON (2)
value SET_ARC_DIRECTION (4102)
value SET_BACKGROUND_COLOR (4103)
value SET_BOUNDS (4109)
value SET_CLIP_BOX (4108)
value SET_FEATURE_IN_REGISTRY (0x00000004)
value SET_FEATURE_ON_PROCESS (0x00000002)
value SET_FEATURE_ON_THREAD (0x00000001)
value SET_FEATURE_ON_THREAD_INTERNET (0x00000040)
value SET_FEATURE_ON_THREAD_INTRANET (0x00000010)
value SET_FEATURE_ON_THREAD_LOCALMACHINE (0x00000008)
value SET_FEATURE_ON_THREAD_RESTRICTED (0x00000080)
value SET_FEATURE_ON_THREAD_TRUSTED (0x00000020)
value SET_MIRROR_MODE (4110)
value SET_POLY_MODE (4104)
value SET_PURGE_FAILURE_MODE_DISABLED (0x00000002)
value SET_PURGE_FAILURE_MODE_ENABLED (0x00000001)
value SET_REPAIR_DISABLED_AND_BUGCHECK_ON_CORRUPT ((0x00000010))
value SET_REPAIR_ENABLED ((0x00000001))
value SET_REPAIR_VALID_MASK ((0x00000019))
value SET_REPAIR_WARN_ABOUT_DATA_LOSS ((0x00000008))
value SET_SCREEN_ANGLE (4105)
value SET_SPREAD (4106)
value SET_TAPE_DRIVE_INFORMATION (1)
value SET_TAPE_MEDIA_INFORMATION (0)
value SEVERITY_ERROR (1)
value SEVERITY_SUCCESS (0)
value SE_ACCESS_CHECK_FLAG_NO_LEARNING_MODE_LOGGING (0x00000008)
value SE_ACCESS_CHECK_VALID_FLAGS (0x00000008)
value SE_DACL_AUTO_INHERITED ((0x0400))
value SE_DACL_AUTO_INHERIT_REQ ((0x0100))
value SE_DACL_DEFAULTED ((0x0008))
value SE_DACL_PRESENT ((0x0004))
value SE_DACL_PROTECTED ((0x1000))
value SE_ERR_ACCESSDENIED (5)
value SE_ERR_ASSOCINCOMPLETE (27)
value SE_ERR_DDEBUSY (30)
value SE_ERR_DDEFAIL (29)
value SE_ERR_DDETIMEOUT (28)
value SE_ERR_DLLNOTFOUND (32)
value SE_ERR_FNF (2)
value SE_ERR_NOASSOC (31)
value SE_ERR_OOM (8)
value SE_ERR_PNF (3)
value SE_ERR_SHARE (26)
value SE_GROUP_DEFAULTED ((0x0002))
value SE_GROUP_ENABLED ((0x00000004L))
value SE_GROUP_ENABLED_BY_DEFAULT ((0x00000002L))
value SE_GROUP_INTEGRITY ((0x00000020L))
value SE_GROUP_INTEGRITY_ENABLED ((0x00000040L))
value SE_GROUP_LOGON_ID ((0xC0000000L))
value SE_GROUP_MANDATORY ((0x00000001L))
value SE_GROUP_OWNER ((0x00000008L))
value SE_GROUP_RESOURCE ((0x20000000L))
value SE_GROUP_USE_FOR_DENY_ONLY ((0x00000010L))
value SE_GROUP_VALID_ATTRIBUTES ((SE_GROUP_MANDATORY | SE_GROUP_ENABLED_BY_DEFAULT | SE_GROUP_ENABLED | SE_GROUP_OWNER | SE_GROUP_USE_FOR_DENY_ONLY | SE_GROUP_LOGON_ID | SE_GROUP_RESOURCE | SE_GROUP_INTEGRITY | SE_GROUP_INTEGRITY_ENABLED))
value SE_OWNER_DEFAULTED ((0x0001))
value SE_PRIVILEGE_ENABLED ((0x00000002L))
value SE_PRIVILEGE_ENABLED_BY_DEFAULT ((0x00000001L))
value SE_PRIVILEGE_REMOVED ((0X00000004L))
value SE_PRIVILEGE_USED_FOR_ACCESS ((0x80000000L))
value SE_PRIVILEGE_VALID_ATTRIBUTES ((SE_PRIVILEGE_ENABLED_BY_DEFAULT | SE_PRIVILEGE_ENABLED | SE_PRIVILEGE_REMOVED | SE_PRIVILEGE_USED_FOR_ACCESS))
value SE_RM_CONTROL_VALID ((0x4000))
value SE_SACL_AUTO_INHERITED ((0x0800))
value SE_SACL_AUTO_INHERIT_REQ ((0x0200))
value SE_SACL_DEFAULTED ((0x0020))
value SE_SACL_PRESENT ((0x0010))
value SE_SACL_PROTECTED ((0x2000))
value SE_SECURITY_DESCRIPTOR_FLAG_NO_ACCESS_FILTER_ACE (0x00000004)
value SE_SECURITY_DESCRIPTOR_FLAG_NO_LABEL_ACE (0x00000002)
value SE_SECURITY_DESCRIPTOR_FLAG_NO_OWNER_ACE (0x00000001)
value SE_SECURITY_DESCRIPTOR_VALID_FLAGS (0x00000007)
value SE_SELF_RELATIVE ((0x8000))
value SE_SIGNING_LEVEL_ANTIMALWARE (SE_SIGNING_LEVEL_CUSTOM_3)
value SE_SIGNING_LEVEL_AUTHENTICODE (0x00000004)
value SE_SIGNING_LEVEL_DEVELOPER (SE_SIGNING_LEVEL_CUSTOM_1)
value SE_SIGNING_LEVEL_DYNAMIC_CODEGEN (0x0000000B)
value SE_SIGNING_LEVEL_ENTERPRISE (0x00000002)
value SE_SIGNING_LEVEL_MICROSOFT (0x00000008)
value SE_SIGNING_LEVEL_STORE (0x00000006)
value SE_SIGNING_LEVEL_UNCHECKED (0x00000000)
value SE_SIGNING_LEVEL_UNSIGNED (0x00000001)
value SE_SIGNING_LEVEL_WINDOWS (0x0000000C)
value SE_SIGNING_LEVEL_WINDOWS_TCB (0x0000000E)
value SG_CONSTRAINED_GROUP (0x02)
value SG_UNCONSTRAINED_GROUP (0x01)
value SHADEBLENDCAPS (120)
value SHAREVISTRING (SHAREVISTRINGA)
value SHDOCAPI (EXTERN_C DECLSPEC_IMPORT HRESULT STDAPICALLTYPE)
value SHERB_NOCONFIRMATION (0x00000001)
value SHERB_NOPROGRESSUI (0x00000002)
value SHERB_NOSOUND (0x00000004)
value SHGFI_ADDOVERLAYS (0x000000020)
value SHGFI_ATTRIBUTES (0x000000800)
value SHGFI_ATTR_SPECIFIED (0x000020000)
value SHGFI_DISPLAYNAME (0x000000200)
value SHGFI_EXETYPE (0x000002000)
value SHGFI_ICON (0x000000100)
value SHGFI_ICONLOCATION (0x000001000)
value SHGFI_LARGEICON (0x000000000)
value SHGFI_LINKOVERLAY (0x000008000)
value SHGFI_OPENICON (0x000000002)
value SHGFI_OVERLAYINDEX (0x000000040)
value SHGFI_PIDL (0x000000008)
value SHGFI_SELECTED (0x000010000)
value SHGFI_SHELLICONSIZE (0x000000004)
value SHGFI_SMALLICON (0x000000001)
value SHGFI_SYSICONINDEX (0x000004000)
value SHGFI_TYPENAME (0x000000400)
value SHGFI_USEFILEATTRIBUTES (0x000000010)
value SHGNLI_NOLNK (0x000000008)
value SHGNLI_NOLOCNAME (0x000000010)
value SHGNLI_NOUNIQUE (0x000000004)
value SHGNLI_PIDL (0x000000001)
value SHGNLI_PREFIXNAME (0x000000002)
value SHGNLI_USEURLEXT (0x000000020)
value SHGSI_ICON (SHGFI_ICON)
value SHGSI_ICONLOCATION (0)
value SHGSI_LARGEICON (SHGFI_LARGEICON)
value SHGSI_LINKOVERLAY (SHGFI_LINKOVERLAY)
value SHGSI_SELECTED (SHGFI_SELECTED)
value SHGSI_SHELLICONSIZE (SHGFI_SHELLICONSIZE)
value SHGSI_SMALLICON (SHGFI_SMALLICON)
value SHGSI_SYSICONINDEX (SHGFI_SYSICONINDEX)
value SHIFTJIS_CHARSET (128)
value SHIFT_PRESSED (0x0010)
value SHIL_EXTRALARGE (2)
value SHIL_JUMBO (4)
value SHIL_LARGE (0)
value SHIL_LAST (SHIL_JUMBO)
value SHIL_SMALL (1)
value SHIL_SYSSMALL (3)
value SHOW_FULLSCREEN (3)
value SHOW_ICONWINDOW (2)
value SHOW_OPENNOACTIVATE (4)
value SHOW_OPENWINDOW (1)
value SHRT_MAX (32767)
value SHRT_MIN ((-32768))
value SHSTDAPI (EXTERN_C DECLSPEC_IMPORT HRESULT STDAPICALLTYPE)
value SHTDN_REASON_FLAG_CLEAN_UI (0x04000000)
value SHTDN_REASON_FLAG_COMMENT_REQUIRED (0x01000000)
value SHTDN_REASON_FLAG_DIRTY_PROBLEM_ID_REQUIRED (0x02000000)
value SHTDN_REASON_FLAG_DIRTY_UI (0x08000000)
value SHTDN_REASON_FLAG_MOBILE_UI_RESERVED (0x10000000)
value SHTDN_REASON_FLAG_PLANNED (0x80000000)
value SHTDN_REASON_FLAG_USER_DEFINED (0x40000000)
value SHTDN_REASON_LEGACY_API ((SHTDN_REASON_MAJOR_LEGACY_API | SHTDN_REASON_FLAG_PLANNED))
value SHTDN_REASON_MAJOR_APPLICATION (0x00040000)
value SHTDN_REASON_MAJOR_HARDWARE (0x00010000)
value SHTDN_REASON_MAJOR_LEGACY_API (0x00070000)
value SHTDN_REASON_MAJOR_NONE (0x00000000)
value SHTDN_REASON_MAJOR_OPERATINGSYSTEM (0x00020000)
value SHTDN_REASON_MAJOR_OTHER (0x00000000)
value SHTDN_REASON_MAJOR_POWER (0x00060000)
value SHTDN_REASON_MAJOR_SOFTWARE (0x00030000)
value SHTDN_REASON_MAJOR_SYSTEM (0x00050000)
value SHTDN_REASON_MINOR_BLUESCREEN (0x0000000F)
value SHTDN_REASON_MINOR_CORDUNPLUGGED (0x0000000b)
value SHTDN_REASON_MINOR_DC_DEMOTION (0x00000022)
value SHTDN_REASON_MINOR_DC_PROMOTION (0x00000021)
value SHTDN_REASON_MINOR_DISK (0x00000007)
value SHTDN_REASON_MINOR_ENVIRONMENT (0x0000000c)
value SHTDN_REASON_MINOR_HARDWARE_DRIVER (0x0000000d)
value SHTDN_REASON_MINOR_HOTFIX (0x00000011)
value SHTDN_REASON_MINOR_HOTFIX_UNINSTALL (0x00000017)
value SHTDN_REASON_MINOR_HUNG (0x00000005)
value SHTDN_REASON_MINOR_INSTALLATION (0x00000002)
value SHTDN_REASON_MINOR_MAINTENANCE (0x00000001)
value SHTDN_REASON_MINOR_MMC (0x00000019)
value SHTDN_REASON_MINOR_NETWORKCARD (0x00000009)
value SHTDN_REASON_MINOR_NETWORK_CONNECTIVITY (0x00000014)
value SHTDN_REASON_MINOR_NONE (0x000000ff)
value SHTDN_REASON_MINOR_OTHER (0x00000000)
value SHTDN_REASON_MINOR_OTHERDRIVER (0x0000000e)
value SHTDN_REASON_MINOR_POWER_SUPPLY (0x0000000a)
value SHTDN_REASON_MINOR_PROCESSOR (0x00000008)
value SHTDN_REASON_MINOR_RECONFIG (0x00000004)
value SHTDN_REASON_MINOR_SECURITY (0x00000013)
value SHTDN_REASON_MINOR_SECURITYFIX (0x00000012)
value SHTDN_REASON_MINOR_SECURITYFIX_UNINSTALL (0x00000018)
value SHTDN_REASON_MINOR_SERVICEPACK (0x00000010)
value SHTDN_REASON_MINOR_SERVICEPACK_UNINSTALL (0x00000016)
value SHTDN_REASON_MINOR_SYSTEMRESTORE (0x0000001a)
value SHTDN_REASON_MINOR_TERMSRV (0x00000020)
value SHTDN_REASON_MINOR_UNSTABLE (0x00000006)
value SHTDN_REASON_MINOR_UPGRADE (0x00000003)
value SHTDN_REASON_MINOR_WMI (0x00000015)
value SHTDN_REASON_UNKNOWN (SHTDN_REASON_MINOR_NONE)
value SHTDN_REASON_VALID_BIT_MASK (0xc0ffffff)
value SHUFFLE_FILE_FLAG_SKIP_INITIALIZING_NEW_CLUSTERS ((0x00000001))
value SHUTDOWN_ARSO (0x00002000)
value SHUTDOWN_CHECK_SAFE_FOR_SERVER (0x00004000)
value SHUTDOWN_FORCE_OTHERS (0x00000001)
value SHUTDOWN_FORCE_SELF (0x00000002)
value SHUTDOWN_GRACE_OVERRIDE (0x00000020)
value SHUTDOWN_HYBRID (0x00000200)
value SHUTDOWN_INSTALL_UPDATES (0x00000040)
value SHUTDOWN_MOBILE_UI (0x00001000)
value SHUTDOWN_NOREBOOT (0x00000010)
value SHUTDOWN_NORETRY (0x00000001)
value SHUTDOWN_POWEROFF (0x00000008)
value SHUTDOWN_RESTART (0x00000004)
value SHUTDOWN_RESTARTAPPS (0x00000080)
value SHUTDOWN_RESTART_BOOTOPTIONS (0x00000400)
value SHUTDOWN_SKIP_SVC_PRESHUTDOWN (0x00000100)
value SHUTDOWN_SOFT_REBOOT (0x00000800)
value SHUTDOWN_SYSTEM_INITIATED (0x00010000)
value SHUTDOWN_TYPE_LEN (32)
value SHUTDOWN_VAIL_CONTAINER (0x00008000)
value SID_HASH_SIZE (32)
value SID_MAX_SUB_AUTHORITIES ((15))
value SID_RECOMMENDED_SUB_AUTHORITIES ((1))
value SID_REVISION ((1))
value SIF_ALL ((SIF_RANGE | SIF_PAGE | SIF_POS | SIF_TRACKPOS))
value SIF_DISABLENOSCROLL (0x0008)
value SIF_PAGE (0x0002)
value SIF_POS (0x0004)
value SIF_RANGE (0x0001)
value SIF_TRACKPOS (0x0010)
value SIID_INVALID (((SHSTOCKICONID)-1))
value SIMPLEBLOB (0x1)
value SIMPLEREGION (2)
value SIMULATED_FONTTYPE (0x8000)
value SITE_PIN_RULES_ALL_SUBDOMAINS_FLAG (0x1)
value SIZEFULLSCREEN (SIZE_MAXIMIZED)
value SIZEICONIC (SIZE_MINIMIZED)
value SIZENORMAL (SIZE_RESTORED)
value SIZEOF_RFPO_DATA (16)
value SIZEPALETTE (104)
value SIZEZOOMHIDE (SIZE_MAXHIDE)
value SIZEZOOMSHOW (SIZE_MAXSHOW)
value SIZE_MAXHIDE (4)
value SIZE_MAXIMIZED (2)
value SIZE_MAXSHOW (3)
value SIZE_MINIMIZED (1)
value SIZE_RESTORED (0)
value SKF_AUDIBLEFEEDBACK (0x00000040)
value SKF_AVAILABLE (0x00000002)
value SKF_CONFIRMHOTKEY (0x00000008)
value SKF_HOTKEYACTIVE (0x00000004)
value SKF_HOTKEYSOUND (0x00000010)
value SKF_INDICATOR (0x00000020)
value SKF_LALTLATCHED (0x10000000)
value SKF_LALTLOCKED (0x00100000)
value SKF_LCTLLATCHED (0x04000000)
value SKF_LCTLLOCKED (0x00040000)
value SKF_LSHIFTLATCHED (0x01000000)
value SKF_LSHIFTLOCKED (0x00010000)
value SKF_LWINLATCHED (0x40000000)
value SKF_LWINLOCKED (0x00400000)
value SKF_RALTLATCHED (0x20000000)
value SKF_RALTLOCKED (0x00200000)
value SKF_RCTLLATCHED (0x08000000)
value SKF_RCTLLOCKED (0x00080000)
value SKF_RSHIFTLATCHED (0x02000000)
value SKF_RSHIFTLOCKED (0x00020000)
value SKF_RWINLATCHED (0x80000000)
value SKF_RWINLOCKED (0x00800000)
value SKF_STICKYKEYSON (0x00000001)
value SKF_TRISTATE (0x00000080)
value SKF_TWOKEYSOFF (0x00000100)
value SLE_ERROR (0x00000001)
value SLE_MINORERROR (0x00000002)
value SLE_WARNING (0x00000003)
value SMART_ABORT_OFFLINE_SELFTEST (127)
value SMART_CMD (0xB0)
value SMART_CYL_HI (0xC2)
value SMART_CYL_LOW (0x4F)
value SMART_ERROR_NO_MEM (7)
value SMART_EXTENDED_SELFTEST_CAPTIVE (130)
value SMART_EXTENDED_SELFTEST_OFFLINE (2)
value SMART_IDE_ERROR (1)
value SMART_INVALID_BUFFER (4)
value SMART_INVALID_COMMAND (3)
value SMART_INVALID_DRIVE (5)
value SMART_INVALID_FLAG (2)
value SMART_INVALID_IOCTL (6)
value SMART_INVALID_REGISTER (8)
value SMART_LOG_SECTOR_SIZE (512)
value SMART_NOT_SUPPORTED (9)
value SMART_NO_ERROR (0)
value SMART_NO_IDE_DEVICE (10)
value SMART_OFFLINE_ROUTINE_OFFLINE (0)
value SMART_READ_LOG (0xD5)
value SMART_SHORT_SELFTEST_CAPTIVE (129)
value SMART_SHORT_SELFTEST_OFFLINE (1)
value SMART_WRITE_LOG (0xd6)
value SMTO_ABORTIFHUNG (0x0002)
value SMTO_BLOCK (0x0001)
value SMTO_ERRORONEXIT (0x0020)
value SMTO_NORMAL (0x0000)
value SMTO_NOTIMEOUTIFNOTHUNG (0x0008)
value SMT_UNPARKING_POLICY_CORE (0)
value SMT_UNPARKING_POLICY_CORE_PER_THREAD (1)
value SMT_UNPARKING_POLICY_LP_ROUNDROBIN (2)
value SMT_UNPARKING_POLICY_LP_SEQUENTIAL (3)
value SM_ARRANGE (56)
value SM_CARETBLINKINGENABLED (0x2002)
value SM_CLEANBOOT (67)
value SM_CMETRICS (97)
value SM_CMONITORS (80)
value SM_CMOUSEBUTTONS (43)
value SM_CONVERTIBLESLATEMODE (0x2003)
value SM_CXBORDER (5)
value SM_CXCURSOR (13)
value SM_CXDLGFRAME (7)
value SM_CXDOUBLECLK (36)
value SM_CXDRAG (68)
value SM_CXEDGE (45)
value SM_CXFIXEDFRAME (SM_CXDLGFRAME)
value SM_CXFOCUSBORDER (83)
value SM_CXFRAME (32)
value SM_CXFULLSCREEN (16)
value SM_CXHSCROLL (21)
value SM_CXHTHUMB (10)
value SM_CXICON (11)
value SM_CXICONSPACING (38)
value SM_CXMAXIMIZED (61)
value SM_CXMAXTRACK (59)
value SM_CXMENUCHECK (71)
value SM_CXMENUSIZE (54)
value SM_CXMIN (28)
value SM_CXMINIMIZED (57)
value SM_CXMINSPACING (47)
value SM_CXMINTRACK (34)
value SM_CXPADDEDBORDER (92)
value SM_CXSCREEN (0)
value SM_CXSIZE (30)
value SM_CXSIZEFRAME (SM_CXFRAME)
value SM_CXSMICON (49)
value SM_CXSMSIZE (52)
value SM_CXVIRTUALSCREEN (78)
value SM_CXVSCROLL (2)
value SM_CYBORDER (6)
value SM_CYCAPTION (4)
value SM_CYCURSOR (14)
value SM_CYDLGFRAME (8)
value SM_CYDOUBLECLK (37)
value SM_CYDRAG (69)
value SM_CYEDGE (46)
value SM_CYFIXEDFRAME (SM_CYDLGFRAME)
value SM_CYFOCUSBORDER (84)
value SM_CYFRAME (33)
value SM_CYFULLSCREEN (17)
value SM_CYHSCROLL (3)
value SM_CYICON (12)
value SM_CYICONSPACING (39)
value SM_CYKANJIWINDOW (18)
value SM_CYMAXIMIZED (62)
value SM_CYMAXTRACK (60)
value SM_CYMENU (15)
value SM_CYMENUCHECK (72)
value SM_CYMENUSIZE (55)
value SM_CYMIN (29)
value SM_CYMINIMIZED (58)
value SM_CYMINSPACING (48)
value SM_CYMINTRACK (35)
value SM_CYSCREEN (1)
value SM_CYSIZE (31)
value SM_CYSIZEFRAME (SM_CYFRAME)
value SM_CYSMCAPTION (51)
value SM_CYSMICON (50)
value SM_CYSMSIZE (53)
value SM_CYVIRTUALSCREEN (79)
value SM_CYVSCROLL (20)
value SM_CYVTHUMB (9)
value SM_DBCSENABLED (42)
value SM_DEBUG (22)
value SM_DIGITIZER (94)
value SM_IMMENABLED (82)
value SM_MAXIMUMTOUCHES (95)
value SM_MEDIACENTER (87)
value SM_MENUDROPALIGNMENT (40)
value SM_MIDEASTENABLED (74)
value SM_MOUSEHORIZONTALWHEELPRESENT (91)
value SM_MOUSEPRESENT (19)
value SM_MOUSEWHEELPRESENT (75)
value SM_NETWORK (63)
value SM_PENWINDOWS (41)
value SM_REMOTECONTROL (0x2001)
value SM_REMOTESESSION (0x1000)
value SM_SAMEDISPLAYFORMAT (81)
value SM_SECURE (44)
value SM_SHOWSOUNDS (70)
value SM_SHUTTINGDOWN (0x2000)
value SM_SLOWMACHINE (73)
value SM_STARTER (88)
value SM_SWAPBUTTON (23)
value SM_SYSTEMDOCKED (0x2004)
value SM_TABLETPC (86)
value SM_XVIRTUALSCREEN (76)
value SM_YVIRTUALSCREEN (77)
value SNAPSHOT_POLICY_ALWAYS (1)
value SNAPSHOT_POLICY_NEVER (0)
value SNAPSHOT_POLICY_UNPLANNED (2)
value SND_ALIAS (0x00010000L)
value SND_ALIAS_ID (0x00110000L)
value SND_ALIAS_START (0)
value SND_APPLICATION (0x0080)
value SND_ASYNC (0x0001)
value SND_FILENAME (0x00020000L)
value SND_LOOP (0x0008)
value SND_MEMORY (0x0004)
value SND_NODEFAULT (0x0002)
value SND_NOSTOP (0x0010)
value SND_NOWAIT (0x00002000L)
value SND_PURGE (0x0040)
value SND_RESOURCE (0x00040004L)
value SND_RING (0x00100000L)
value SND_SENTRY (0x00080000L)
value SND_SYNC (0x0000)
value SND_SYSTEM (0x00200000L)
value SOCKET_ERROR ((-1))
value SOCK_DGRAM (2)
value SOCK_NOTIFY_EVENTS_ALL ((SOCK_NOTIFY_REGISTER_EVENTS_ALL | SOCK_NOTIFY_EVENT_ERR | SOCK_NOTIFY_EVENT_REMOVE))
value SOCK_NOTIFY_EVENT_ERR (0x40)
value SOCK_NOTIFY_EVENT_HANGUP (SOCK_NOTIFY_REGISTER_EVENT_HANGUP)
value SOCK_NOTIFY_EVENT_IN (SOCK_NOTIFY_REGISTER_EVENT_IN)
value SOCK_NOTIFY_EVENT_OUT (SOCK_NOTIFY_REGISTER_EVENT_OUT)
value SOCK_NOTIFY_EVENT_REMOVE (0x80)
value SOCK_NOTIFY_OP_DISABLE (0x02)
value SOCK_NOTIFY_OP_ENABLE (0x01)
value SOCK_NOTIFY_OP_NONE (0x00)
value SOCK_NOTIFY_OP_REMOVE (0x04)
value SOCK_NOTIFY_REGISTER_EVENTS_ALL ((SOCK_NOTIFY_REGISTER_EVENT_IN | SOCK_NOTIFY_REGISTER_EVENT_OUT | SOCK_NOTIFY_REGISTER_EVENT_HANGUP))
value SOCK_NOTIFY_REGISTER_EVENT_HANGUP (0x04)
value SOCK_NOTIFY_REGISTER_EVENT_IN (0x01)
value SOCK_NOTIFY_REGISTER_EVENT_NONE (0x00)
value SOCK_NOTIFY_REGISTER_EVENT_OUT (0x02)
value SOCK_NOTIFY_TRIGGER_ALL ((SOCK_NOTIFY_TRIGGER_ONESHOT | SOCK_NOTIFY_TRIGGER_PERSISTENT | SOCK_NOTIFY_TRIGGER_LEVEL | SOCK_NOTIFY_TRIGGER_EDGE))
value SOCK_NOTIFY_TRIGGER_EDGE (0x08)
value SOCK_NOTIFY_TRIGGER_LEVEL (0x04)
value SOCK_NOTIFY_TRIGGER_ONESHOT (0x01)
value SOCK_NOTIFY_TRIGGER_PERSISTENT (0x02)
value SOCK_RAW (3)
value SOCK_RDM (4)
value SOCK_SEQPACKET (5)
value SOCK_STREAM (1)
value SOFTDIST_ADSTATE_AVAILABLE (0x00000001)
value SOFTDIST_ADSTATE_DOWNLOADED (0x00000002)
value SOFTDIST_ADSTATE_INSTALLED (0x00000003)
value SOFTDIST_ADSTATE_NONE (0x00000000)
value SOFTDIST_FLAG_DELETE_SUBSCRIPTION (0x00000008)
value SOFTDIST_FLAG_USAGE_AUTOINSTALL (0x00000004)
value SOFTDIST_FLAG_USAGE_EMAIL (0x00000001)
value SOFTDIST_FLAG_USAGE_PRECACHE (0x00000002)
value SOL_IP ((SOL_SOCKET-4))
value SOL_SOCKET (0xffff)
value SOMAXCONN (0x7fffffff)
value SORTED_CTL_EXT_HASHED_SUBJECT_IDENTIFIER_FLAG (0x1)
value SORTING_PARADIGM_ICU (0x01000000)
value SORTING_PARADIGM_NLS (0x00000000)
value SORT_CHINESE_BOPOMOFO (0x3)
value SORT_CHINESE_PRC (0x2)
value SORT_CHINESE_PRCP (0x0)
value SORT_CHINESE_RADICALSTROKE (0x4)
value SORT_CHINESE_UNICODE (0x1)
value SORT_DEFAULT (0x0)
value SORT_DIGITSASNUMBERS (0x00000008)
value SORT_GEORGIAN_MODERN (0x1)
value SORT_GEORGIAN_TRADITIONAL (0x0)
value SORT_GERMAN_PHONE_BOOK (0x1)
value SORT_HUNGARIAN_DEFAULT (0x0)
value SORT_HUNGARIAN_TECHNICAL (0x1)
value SORT_INVARIANT_MATH (0x1)
value SORT_JAPANESE_RADICALSTROKE (0x4)
value SORT_JAPANESE_UNICODE (0x1)
value SORT_JAPANESE_XJIS (0x0)
value SORT_KOREAN_KSC (0x0)
value SORT_KOREAN_UNICODE (0x1)
value SORT_STRINGSORT (0x00001000)
value SOUND_SYSTEM_APPEND (14)
value SOUND_SYSTEM_APPSTART (12)
value SOUND_SYSTEM_BEEP (3)
value SOUND_SYSTEM_ERROR (4)
value SOUND_SYSTEM_FAULT (13)
value SOUND_SYSTEM_INFORMATION (7)
value SOUND_SYSTEM_MAXIMIZE (8)
value SOUND_SYSTEM_MENUCOMMAND (15)
value SOUND_SYSTEM_MENUPOPUP (16)
value SOUND_SYSTEM_MINIMIZE (9)
value SOUND_SYSTEM_QUESTION (5)
value SOUND_SYSTEM_RESTOREDOWN (11)
value SOUND_SYSTEM_RESTOREUP (10)
value SOUND_SYSTEM_SHUTDOWN (2)
value SOUND_SYSTEM_STARTUP (1)
value SOUND_SYSTEM_WARNING (6)
value SO_ACCEPTCONN (0x0002)
value SO_BROADCAST (0x0020)
value SO_BSP_STATE (0x1009)
value SO_COMPARTMENT_ID (0x3004)
value SO_CONDITIONAL_ACCEPT (0x3002)
value SO_DEBUG (0x0001)
value SO_DONTROUTE (0x0010)
value SO_ERROR (0x1007)
value SO_GROUP_ID (0x2001)
value SO_GROUP_PRIORITY (0x2002)
value SO_KEEPALIVE (0x0008)
value SO_LINGER (0x0080)
value SO_MAX_MSG_SIZE (0x2003)
value SO_OOBINLINE (0x0100)
value SO_ORIGINAL_DST (0x300F)
value SO_PAUSE_ACCEPT (0x3003)
value SO_PORT_SCALABILITY (0x3006)
value SO_PROTOCOL_INFO (SO_PROTOCOL_INFOA)
value SO_PROTOCOL_INFOA (0x2004)
value SO_PROTOCOL_INFOW (0x2005)
value SO_RANDOMIZE_PORT (0x3005)
value SO_RCVBUF (0x1002)
value SO_RCVLOWAT (0x1004)
value SO_RCVTIMEO (0x1006)
value SO_REUSEADDR (0x0004)
value SO_REUSE_MULTICASTPORT (0x3008)
value SO_REUSE_UNICASTPORT (0x3007)
value SO_SNDBUF (0x1001)
value SO_SNDLOWAT (0x1003)
value SO_SNDTIMEO (0x1005)
value SO_TYPE (0x1008)
value SO_USELOOPBACK (0x0040)
value SPACEPARITY (4)
value SPACES_TRACKED_OFFSET_HEADER_FLAG (0x0002)
value SPAPI_E_AUTHENTICODE_DISALLOWED (_HRESULT_TYPEDEF_(0x800F0240L))
value SPAPI_E_AUTHENTICODE_PUBLISHER_NOT_TRUSTED (_HRESULT_TYPEDEF_(0x800F0243L))
value SPAPI_E_AUTHENTICODE_TRUSTED_PUBLISHER (_HRESULT_TYPEDEF_(0x800F0241L))
value SPAPI_E_AUTHENTICODE_TRUST_NOT_ESTABLISHED (_HRESULT_TYPEDEF_(0x800F0242L))
value SPAPI_E_BAD_INTERFACE_INSTALLSECT (_HRESULT_TYPEDEF_(0x800F021DL))
value SPAPI_E_BAD_SECTION_NAME_LINE (_HRESULT_TYPEDEF_(0x800F0001L))
value SPAPI_E_BAD_SERVICE_INSTALLSECT (_HRESULT_TYPEDEF_(0x800F0217L))
value SPAPI_E_CANT_LOAD_CLASS_ICON (_HRESULT_TYPEDEF_(0x800F020CL))
value SPAPI_E_CANT_REMOVE_DEVINST (_HRESULT_TYPEDEF_(0x800F0232L))
value SPAPI_E_CLASS_MISMATCH (_HRESULT_TYPEDEF_(0x800F0201L))
value SPAPI_E_DEVICE_INSTALLER_NOT_READY (_HRESULT_TYPEDEF_(0x800F0246L))
value SPAPI_E_DEVICE_INSTALL_BLOCKED (_HRESULT_TYPEDEF_(0x800F0248L))
value SPAPI_E_DEVICE_INTERFACE_ACTIVE (_HRESULT_TYPEDEF_(0x800F021BL))
value SPAPI_E_DEVICE_INTERFACE_REMOVED (_HRESULT_TYPEDEF_(0x800F021CL))
value SPAPI_E_DEVINFO_DATA_LOCKED (_HRESULT_TYPEDEF_(0x800F0213L))
value SPAPI_E_DEVINFO_LIST_LOCKED (_HRESULT_TYPEDEF_(0x800F0212L))
value SPAPI_E_DEVINFO_NOT_REGISTERED (_HRESULT_TYPEDEF_(0x800F0208L))
value SPAPI_E_DEVINSTALL_QUEUE_NONNATIVE (_HRESULT_TYPEDEF_(0x800F0230L))
value SPAPI_E_DEVINST_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x800F0207L))
value SPAPI_E_DI_BAD_PATH (_HRESULT_TYPEDEF_(0x800F0214L))
value SPAPI_E_DI_DONT_INSTALL (_HRESULT_TYPEDEF_(0x800F022BL))
value SPAPI_E_DI_DO_DEFAULT (_HRESULT_TYPEDEF_(0x800F020EL))
value SPAPI_E_DI_FUNCTION_OBSOLETE (_HRESULT_TYPEDEF_(0x800F023EL))
value SPAPI_E_DI_NOFILECOPY (_HRESULT_TYPEDEF_(0x800F020FL))
value SPAPI_E_DI_POSTPROCESSING_REQUIRED (_HRESULT_TYPEDEF_(0x800F0226L))
value SPAPI_E_DRIVER_INSTALL_BLOCKED (_HRESULT_TYPEDEF_(0x800F0249L))
value SPAPI_E_DRIVER_NONNATIVE (_HRESULT_TYPEDEF_(0x800F0234L))
value SPAPI_E_DRIVER_STORE_ADD_FAILED (_HRESULT_TYPEDEF_(0x800F0247L))
value SPAPI_E_DRIVER_STORE_DELETE_FAILED (_HRESULT_TYPEDEF_(0x800F024CL))
value SPAPI_E_DUPLICATE_FOUND (_HRESULT_TYPEDEF_(0x800F0202L))
value SPAPI_E_ERROR_NOT_INSTALLED (_HRESULT_TYPEDEF_(0x800F1000L))
value SPAPI_E_EXPECTED_SECTION_NAME (_HRESULT_TYPEDEF_(0x800F0000L))
value SPAPI_E_FILEQUEUE_LOCKED (_HRESULT_TYPEDEF_(0x800F0216L))
value SPAPI_E_FILE_HASH_NOT_IN_CATALOG (_HRESULT_TYPEDEF_(0x800F024BL))
value SPAPI_E_GENERAL_SYNTAX (_HRESULT_TYPEDEF_(0x800F0003L))
value SPAPI_E_INCORRECTLY_COPIED_INF (_HRESULT_TYPEDEF_(0x800F0237L))
value SPAPI_E_INF_IN_USE_BY_DEVICES (_HRESULT_TYPEDEF_(0x800F023DL))
value SPAPI_E_INVALID_CLASS (_HRESULT_TYPEDEF_(0x800F0206L))
value SPAPI_E_INVALID_CLASS_INSTALLER (_HRESULT_TYPEDEF_(0x800F020DL))
value SPAPI_E_INVALID_COINSTALLER (_HRESULT_TYPEDEF_(0x800F0227L))
value SPAPI_E_INVALID_DEVINST_NAME (_HRESULT_TYPEDEF_(0x800F0205L))
value SPAPI_E_INVALID_FILTER_DRIVER (_HRESULT_TYPEDEF_(0x800F022CL))
value SPAPI_E_INVALID_HWPROFILE (_HRESULT_TYPEDEF_(0x800F0210L))
value SPAPI_E_INVALID_INF_LOGCONFIG (_HRESULT_TYPEDEF_(0x800F022AL))
value SPAPI_E_INVALID_MACHINENAME (_HRESULT_TYPEDEF_(0x800F0220L))
value SPAPI_E_INVALID_PROPPAGE_PROVIDER (_HRESULT_TYPEDEF_(0x800F0224L))
value SPAPI_E_INVALID_REFERENCE_STRING (_HRESULT_TYPEDEF_(0x800F021FL))
value SPAPI_E_INVALID_REG_PROPERTY (_HRESULT_TYPEDEF_(0x800F0209L))
value SPAPI_E_INVALID_TARGET (_HRESULT_TYPEDEF_(0x800F0233L))
value SPAPI_E_KEY_DOES_NOT_EXIST (_HRESULT_TYPEDEF_(0x800F0204L))
value SPAPI_E_LINE_NOT_FOUND (_HRESULT_TYPEDEF_(0x800F0102L))
value SPAPI_E_MACHINE_UNAVAILABLE (_HRESULT_TYPEDEF_(0x800F0222L))
value SPAPI_E_NON_WINDOWS_DRIVER (_HRESULT_TYPEDEF_(0x800F022EL))
value SPAPI_E_NON_WINDOWS_NT_DRIVER (_HRESULT_TYPEDEF_(0x800F022DL))
value SPAPI_E_NOT_AN_INSTALLED_OEM_INF (_HRESULT_TYPEDEF_(0x800F023CL))
value SPAPI_E_NOT_DISABLEABLE (_HRESULT_TYPEDEF_(0x800F0231L))
value SPAPI_E_NO_ASSOCIATED_CLASS (_HRESULT_TYPEDEF_(0x800F0200L))
value SPAPI_E_NO_ASSOCIATED_SERVICE (_HRESULT_TYPEDEF_(0x800F0219L))
value SPAPI_E_NO_AUTHENTICODE_CATALOG (_HRESULT_TYPEDEF_(0x800F023FL))
value SPAPI_E_NO_BACKUP (_HRESULT_TYPEDEF_(0x800F0103L))
value SPAPI_E_NO_CATALOG_FOR_OEM_INF (_HRESULT_TYPEDEF_(0x800F022FL))
value SPAPI_E_NO_CLASSINSTALL_PARAMS (_HRESULT_TYPEDEF_(0x800F0215L))
value SPAPI_E_NO_CLASS_DRIVER_LIST (_HRESULT_TYPEDEF_(0x800F0218L))
value SPAPI_E_NO_COMPAT_DRIVERS (_HRESULT_TYPEDEF_(0x800F0228L))
value SPAPI_E_NO_CONFIGMGR_SERVICES (_HRESULT_TYPEDEF_(0x800F0223L))
value SPAPI_E_NO_DEFAULT_DEVICE_INTERFACE (_HRESULT_TYPEDEF_(0x800F021AL))
value SPAPI_E_NO_DEVICE_ICON (_HRESULT_TYPEDEF_(0x800F0229L))
value SPAPI_E_NO_DEVICE_SELECTED (_HRESULT_TYPEDEF_(0x800F0211L))
value SPAPI_E_NO_DRIVER_SELECTED (_HRESULT_TYPEDEF_(0x800F0203L))
value SPAPI_E_NO_INF (_HRESULT_TYPEDEF_(0x800F020AL))
value SPAPI_E_NO_SUCH_DEVICE_INTERFACE (_HRESULT_TYPEDEF_(0x800F0225L))
value SPAPI_E_NO_SUCH_DEVINST (_HRESULT_TYPEDEF_(0x800F020BL))
value SPAPI_E_NO_SUCH_INTERFACE_CLASS (_HRESULT_TYPEDEF_(0x800F021EL))
value SPAPI_E_ONLY_VALIDATE_VIA_AUTHENTICODE (_HRESULT_TYPEDEF_(0x800F0245L))
value SPAPI_E_PNP_REGISTRY_ERROR (_HRESULT_TYPEDEF_(0x800F023AL))
value SPAPI_E_REMOTE_COMM_FAILURE (_HRESULT_TYPEDEF_(0x800F0221L))
value SPAPI_E_REMOTE_REQUEST_UNSUPPORTED (_HRESULT_TYPEDEF_(0x800F023BL))
value SPAPI_E_SCE_DISABLED (_HRESULT_TYPEDEF_(0x800F0238L))
value SPAPI_E_SECTION_NAME_TOO_LONG (_HRESULT_TYPEDEF_(0x800F0002L))
value SPAPI_E_SECTION_NOT_FOUND (_HRESULT_TYPEDEF_(0x800F0101L))
value SPAPI_E_SET_SYSTEM_RESTORE_POINT (_HRESULT_TYPEDEF_(0x800F0236L))
value SPAPI_E_SIGNATURE_OSATTRIBUTE_MISMATCH (_HRESULT_TYPEDEF_(0x800F0244L))
value SPAPI_E_UNKNOWN_EXCEPTION (_HRESULT_TYPEDEF_(0x800F0239L))
value SPAPI_E_UNRECOVERABLE_STACK_OVERFLOW (_HRESULT_TYPEDEF_(0x800F0300L))
value SPAPI_E_WRONG_INF_STYLE (_HRESULT_TYPEDEF_(0x800F0100L))
value SPAPI_E_WRONG_INF_TYPE (_HRESULT_TYPEDEF_(0x800F024AL))
value SPECIFIC_RIGHTS_ALL ((0x0000FFFFL))
value SPIF_SENDCHANGE (SPIF_SENDWININICHANGE)
value SPIF_SENDWININICHANGE (0x0002)
value SPIF_UPDATEINIFILE (0x0001)
value SPI_GETACCESSTIMEOUT (0x003C)
value SPI_GETACTIVEWINDOWTRACKING (0x1000)
value SPI_GETACTIVEWNDTRKTIMEOUT (0x2002)
value SPI_GETACTIVEWNDTRKZORDER (0x100C)
value SPI_GETANIMATION (0x0048)
value SPI_GETAUDIODESCRIPTION (0x0074)
value SPI_GETBEEP (0x0001)
value SPI_GETBLOCKSENDINPUTRESETS (0x1026)
value SPI_GETBORDER (0x0005)
value SPI_GETCARETBROWSING (0x104C)
value SPI_GETCARETTIMEOUT (0x2022)
value SPI_GETCARETWIDTH (0x2006)
value SPI_GETCLEARTYPE (0x1048)
value SPI_GETCLIENTAREAANIMATION (0x1042)
value SPI_GETCOMBOBOXANIMATION (0x1004)
value SPI_GETCONTACTVISUALIZATION (0x2018)
value SPI_GETCURSORSHADOW (0x101A)
value SPI_GETDEFAULTINPUTLANG (0x0059)
value SPI_GETDESKWALLPAPER (0x0073)
value SPI_GETDISABLEOVERLAPPEDCONTENT (0x1040)
value SPI_GETDOCKMOVING (0x0090)
value SPI_GETDRAGFROMMAXIMIZE (0x008C)
value SPI_GETDRAGFULLWINDOWS (0x0026)
value SPI_GETDROPSHADOW (0x1024)
value SPI_GETFASTTASKSWITCH (0x0023)
value SPI_GETFILTERKEYS (0x0032)
value SPI_GETFLATMENU (0x1022)
value SPI_GETFOCUSBORDERHEIGHT (0x2010)
value SPI_GETFOCUSBORDERWIDTH (0x200E)
value SPI_GETFONTSMOOTHING (0x004A)
value SPI_GETFONTSMOOTHINGCONTRAST (0x200C)
value SPI_GETFONTSMOOTHINGORIENTATION (0x2012)
value SPI_GETFONTSMOOTHINGTYPE (0x200A)
value SPI_GETFOREGROUNDFLASHCOUNT (0x2004)
value SPI_GETFOREGROUNDLOCKTIMEOUT (0x2000)
value SPI_GETGESTUREVISUALIZATION (0x201A)
value SPI_GETGRADIENTCAPTIONS (0x1008)
value SPI_GETGRIDGRANULARITY (0x0012)
value SPI_GETHANDEDNESS (0x2024)
value SPI_GETHIGHCONTRAST (0x0042)
value SPI_GETHOTTRACKING (0x100E)
value SPI_GETHUNGAPPTIMEOUT (0x0078)
value SPI_GETICONMETRICS (0x002D)
value SPI_GETICONTITLELOGFONT (0x001F)
value SPI_GETICONTITLEWRAP (0x0019)
value SPI_GETKEYBOARDCUES (0x100A)
value SPI_GETKEYBOARDDELAY (0x0016)
value SPI_GETKEYBOARDPREF (0x0044)
value SPI_GETKEYBOARDSPEED (0x000A)
value SPI_GETLISTBOXSMOOTHSCROLLING (0x1006)
value SPI_GETLOGICALDPIOVERRIDE (0x009E)
value SPI_GETLOWPOWERACTIVE (0x0053)
value SPI_GETLOWPOWERTIMEOUT (0x004F)
value SPI_GETMENUANIMATION (0x1002)
value SPI_GETMENUDROPALIGNMENT (0x001B)
value SPI_GETMENUFADE (0x1012)
value SPI_GETMENURECT (0x00A2)
value SPI_GETMENUSHOWDELAY (0x006A)
value SPI_GETMENUUNDERLINES (SPI_GETKEYBOARDCUES)
value SPI_GETMESSAGEDURATION (0x2016)
value SPI_GETMINIMIZEDMETRICS (0x002B)
value SPI_GETMINIMUMHITRADIUS (0x2014)
value SPI_GETMOUSE (0x0003)
value SPI_GETMOUSECLICKLOCK (0x101E)
value SPI_GETMOUSECLICKLOCKTIME (0x2008)
value SPI_GETMOUSEDOCKTHRESHOLD (0x007E)
value SPI_GETMOUSEDRAGOUTTHRESHOLD (0x0084)
value SPI_GETMOUSEHOVERHEIGHT (0x0064)
value SPI_GETMOUSEHOVERTIME (0x0066)
value SPI_GETMOUSEHOVERWIDTH (0x0062)
value SPI_GETMOUSEKEYS (0x0036)
value SPI_GETMOUSESIDEMOVETHRESHOLD (0x0088)
value SPI_GETMOUSESONAR (0x101C)
value SPI_GETMOUSESPEED (0x0070)
value SPI_GETMOUSETRAILS (0x005E)
value SPI_GETMOUSEVANISH (0x1020)
value SPI_GETMOUSEWHEELROUTING (0x201C)
value SPI_GETNONCLIENTMETRICS (0x0029)
value SPI_GETPENARBITRATIONTYPE (0x2020)
value SPI_GETPENDOCKTHRESHOLD (0x0080)
value SPI_GETPENDRAGOUTTHRESHOLD (0x0086)
value SPI_GETPENSIDEMOVETHRESHOLD (0x008A)
value SPI_GETPENVISUALIZATION (0x201E)
value SPI_GETPOWEROFFACTIVE (0x0054)
value SPI_GETPOWEROFFTIMEOUT (0x0050)
value SPI_GETSCREENREADER (0x0046)
value SPI_GETSCREENSAVEACTIVE (0x0010)
value SPI_GETSCREENSAVERRUNNING (0x0072)
value SPI_GETSCREENSAVESECURE (0x0076)
value SPI_GETSCREENSAVETIMEOUT (0x000E)
value SPI_GETSELECTIONFADE (0x1014)
value SPI_GETSERIALKEYS (0x003E)
value SPI_GETSHOWIMEUI (0x006E)
value SPI_GETSHOWSOUNDS (0x0038)
value SPI_GETSNAPSIZING (0x008E)
value SPI_GETSNAPTODEFBUTTON (0x005F)
value SPI_GETSOUNDSENTRY (0x0040)
value SPI_GETSPEECHRECOGNITION (0x104A)
value SPI_GETSTICKYKEYS (0x003A)
value SPI_GETSYSTEMLANGUAGEBAR (0x1050)
value SPI_GETTHREADLOCALINPUTSETTINGS (0x104E)
value SPI_GETTOGGLEKEYS (0x0034)
value SPI_GETTOOLTIPANIMATION (0x1016)
value SPI_GETTOOLTIPFADE (0x1018)
value SPI_GETTOUCHPREDICTIONPARAMETERS (0x009C)
value SPI_GETUIEFFECTS (0x103E)
value SPI_GETWAITTOKILLSERVICETIMEOUT (0x007C)
value SPI_GETWAITTOKILLTIMEOUT (0x007A)
value SPI_GETWHEELSCROLLCHARS (0x006C)
value SPI_GETWHEELSCROLLLINES (0x0068)
value SPI_GETWINARRANGING (0x0082)
value SPI_GETWINDOWSEXTENSION (0x005C)
value SPI_GETWORKAREA (0x0030)
value SPI_ICONHORIZONTALSPACING (0x000D)
value SPI_ICONVERTICALSPACING (0x0018)
value SPI_LANGDRIVER (0x000C)
value SPI_SCREENSAVERRUNNING (SPI_SETSCREENSAVERRUNNING)
value SPI_SETACCESSTIMEOUT (0x003D)
value SPI_SETACTIVEWINDOWTRACKING (0x1001)
value SPI_SETACTIVEWNDTRKTIMEOUT (0x2003)
value SPI_SETACTIVEWNDTRKZORDER (0x100D)
value SPI_SETANIMATION (0x0049)
value SPI_SETAUDIODESCRIPTION (0x0075)
value SPI_SETBEEP (0x0002)
value SPI_SETBLOCKSENDINPUTRESETS (0x1027)
value SPI_SETBORDER (0x0006)
value SPI_SETCARETBROWSING (0x104D)
value SPI_SETCARETTIMEOUT (0x2023)
value SPI_SETCARETWIDTH (0x2007)
value SPI_SETCLEARTYPE (0x1049)
value SPI_SETCLIENTAREAANIMATION (0x1043)
value SPI_SETCOMBOBOXANIMATION (0x1005)
value SPI_SETCONTACTVISUALIZATION (0x2019)
value SPI_SETCURSORS (0x0057)
value SPI_SETCURSORSHADOW (0x101B)
value SPI_SETDEFAULTINPUTLANG (0x005A)
value SPI_SETDESKPATTERN (0x0015)
value SPI_SETDESKWALLPAPER (0x0014)
value SPI_SETDISABLEOVERLAPPEDCONTENT (0x1041)
value SPI_SETDOCKMOVING (0x0091)
value SPI_SETDOUBLECLICKTIME (0x0020)
value SPI_SETDOUBLECLKHEIGHT (0x001E)
value SPI_SETDOUBLECLKWIDTH (0x001D)
value SPI_SETDRAGFROMMAXIMIZE (0x008D)
value SPI_SETDRAGFULLWINDOWS (0x0025)
value SPI_SETDRAGHEIGHT (0x004D)
value SPI_SETDRAGWIDTH (0x004C)
value SPI_SETDROPSHADOW (0x1025)
value SPI_SETFASTTASKSWITCH (0x0024)
value SPI_SETFILTERKEYS (0x0033)
value SPI_SETFLATMENU (0x1023)
value SPI_SETFOCUSBORDERHEIGHT (0x2011)
value SPI_SETFOCUSBORDERWIDTH (0x200F)
value SPI_SETFONTSMOOTHING (0x004B)
value SPI_SETFONTSMOOTHINGCONTRAST (0x200D)
value SPI_SETFONTSMOOTHINGORIENTATION (0x2013)
value SPI_SETFONTSMOOTHINGTYPE (0x200B)
value SPI_SETFOREGROUNDFLASHCOUNT (0x2005)
value SPI_SETFOREGROUNDLOCKTIMEOUT (0x2001)
value SPI_SETGESTUREVISUALIZATION (0x201B)
value SPI_SETGRADIENTCAPTIONS (0x1009)
value SPI_SETGRIDGRANULARITY (0x0013)
value SPI_SETHANDEDNESS (0x2025)
value SPI_SETHANDHELD (0x004E)
value SPI_SETHIGHCONTRAST (0x0043)
value SPI_SETHOTTRACKING (0x100F)
value SPI_SETHUNGAPPTIMEOUT (0x0079)
value SPI_SETICONMETRICS (0x002E)
value SPI_SETICONS (0x0058)
value SPI_SETICONTITLELOGFONT (0x0022)
value SPI_SETICONTITLEWRAP (0x001A)
value SPI_SETKEYBOARDCUES (0x100B)
value SPI_SETKEYBOARDDELAY (0x0017)
value SPI_SETKEYBOARDPREF (0x0045)
value SPI_SETKEYBOARDSPEED (0x000B)
value SPI_SETLANGTOGGLE (0x005B)
value SPI_SETLISTBOXSMOOTHSCROLLING (0x1007)
value SPI_SETLOGICALDPIOVERRIDE (0x009F)
value SPI_SETLOWPOWERACTIVE (0x0055)
value SPI_SETLOWPOWERTIMEOUT (0x0051)
value SPI_SETMENUANIMATION (0x1003)
value SPI_SETMENUDROPALIGNMENT (0x001C)
value SPI_SETMENUFADE (0x1013)
value SPI_SETMENURECT (0x00A3)
value SPI_SETMENUSHOWDELAY (0x006B)
value SPI_SETMENUUNDERLINES (SPI_SETKEYBOARDCUES)
value SPI_SETMESSAGEDURATION (0x2017)
value SPI_SETMINIMIZEDMETRICS (0x002C)
value SPI_SETMINIMUMHITRADIUS (0x2015)
value SPI_SETMOUSE (0x0004)
value SPI_SETMOUSEBUTTONSWAP (0x0021)
value SPI_SETMOUSECLICKLOCK (0x101F)
value SPI_SETMOUSECLICKLOCKTIME (0x2009)
value SPI_SETMOUSEDOCKTHRESHOLD (0x007F)
value SPI_SETMOUSEDRAGOUTTHRESHOLD (0x0085)
value SPI_SETMOUSEHOVERHEIGHT (0x0065)
value SPI_SETMOUSEHOVERTIME (0x0067)
value SPI_SETMOUSEHOVERWIDTH (0x0063)
value SPI_SETMOUSEKEYS (0x0037)
value SPI_SETMOUSESIDEMOVETHRESHOLD (0x0089)
value SPI_SETMOUSESONAR (0x101D)
value SPI_SETMOUSESPEED (0x0071)
value SPI_SETMOUSETRAILS (0x005D)
value SPI_SETMOUSEVANISH (0x1021)
value SPI_SETMOUSEWHEELROUTING (0x201D)
value SPI_SETNONCLIENTMETRICS (0x002A)
value SPI_SETPENARBITRATIONTYPE (0x2021)
value SPI_SETPENDOCKTHRESHOLD (0x0081)
value SPI_SETPENDRAGOUTTHRESHOLD (0x0087)
value SPI_SETPENSIDEMOVETHRESHOLD (0x008B)
value SPI_SETPENVISUALIZATION (0x201F)
value SPI_SETPENWINDOWS (0x0031)
value SPI_SETPOWEROFFACTIVE (0x0056)
value SPI_SETPOWEROFFTIMEOUT (0x0052)
value SPI_SETSCREENREADER (0x0047)
value SPI_SETSCREENSAVEACTIVE (0x0011)
value SPI_SETSCREENSAVERRUNNING (0x0061)
value SPI_SETSCREENSAVESECURE (0x0077)
value SPI_SETSCREENSAVETIMEOUT (0x000F)
value SPI_SETSELECTIONFADE (0x1015)
value SPI_SETSERIALKEYS (0x003F)
value SPI_SETSHOWIMEUI (0x006F)
value SPI_SETSHOWSOUNDS (0x0039)
value SPI_SETSNAPSIZING (0x008F)
value SPI_SETSNAPTODEFBUTTON (0x0060)
value SPI_SETSOUNDSENTRY (0x0041)
value SPI_SETSPEECHRECOGNITION (0x104B)
value SPI_SETSTICKYKEYS (0x003B)
value SPI_SETSYSTEMLANGUAGEBAR (0x1051)
value SPI_SETTHREADLOCALINPUTSETTINGS (0x104F)
value SPI_SETTOGGLEKEYS (0x0035)
value SPI_SETTOOLTIPANIMATION (0x1017)
value SPI_SETTOOLTIPFADE (0x1019)
value SPI_SETTOUCHPREDICTIONPARAMETERS (0x009D)
value SPI_SETUIEFFECTS (0x103F)
value SPI_SETWAITTOKILLSERVICETIMEOUT (0x007D)
value SPI_SETWAITTOKILLTIMEOUT (0x007B)
value SPI_SETWHEELSCROLLCHARS (0x006D)
value SPI_SETWHEELSCROLLLINES (0x0069)
value SPI_SETWINARRANGING (0x0083)
value SPI_SETWORKAREA (0x002F)
value SPOOL_FILE_PERSISTENT (0x00000001)
value SPOOL_FILE_TEMPORARY (0x00000002)
value SPVERSION_MASK (0x0000FF00)
value SP_APPABORT ((-2))
value SP_BAUD (((DWORD)0x0002))
value SP_DATABITS (((DWORD)0x0004))
value SP_ERROR ((-1))
value SP_HANDSHAKING (((DWORD)0x0010))
value SP_NOTREPORTED (0x4000)
value SP_OUTOFDISK ((-4))
value SP_OUTOFMEMORY ((-5))
value SP_PARITY (((DWORD)0x0001))
value SP_PARITY_CHECK (((DWORD)0x0020))
value SP_RLSD (((DWORD)0x0040))
value SP_SERIALCOMM (((DWORD)0x00000001))
value SP_STOPBITS (((DWORD)0x0008))
value SP_USERABORT ((-3))
value SQLITE_E_ABORT (_HRESULT_TYPEDEF_(0x87AF0004L))
value SQLITE_E_ABORT_ROLLBACK (_HRESULT_TYPEDEF_(0x87AF0204L))
value SQLITE_E_AUTH (_HRESULT_TYPEDEF_(0x87AF0017L))
value SQLITE_E_BUSY (_HRESULT_TYPEDEF_(0x87AF0005L))
value SQLITE_E_BUSY_RECOVERY (_HRESULT_TYPEDEF_(0x87AF0105L))
value SQLITE_E_BUSY_SNAPSHOT (_HRESULT_TYPEDEF_(0x87AF0205L))
value SQLITE_E_CANTOPEN (_HRESULT_TYPEDEF_(0x87AF000EL))
value SQLITE_E_CANTOPEN_CONVPATH (_HRESULT_TYPEDEF_(0x87AF040EL))
value SQLITE_E_CANTOPEN_FULLPATH (_HRESULT_TYPEDEF_(0x87AF030EL))
value SQLITE_E_CANTOPEN_ISDIR (_HRESULT_TYPEDEF_(0x87AF020EL))
value SQLITE_E_CANTOPEN_NOTEMPDIR (_HRESULT_TYPEDEF_(0x87AF010EL))
value SQLITE_E_CONSTRAINT (_HRESULT_TYPEDEF_(0x87AF0013L))
value SQLITE_E_CONSTRAINT_CHECK (_HRESULT_TYPEDEF_(0x87AF0113L))
value SQLITE_E_CONSTRAINT_COMMITHOOK (_HRESULT_TYPEDEF_(0x87AF0213L))
value SQLITE_E_CONSTRAINT_FOREIGNKEY (_HRESULT_TYPEDEF_(0x87AF0313L))
value SQLITE_E_CONSTRAINT_FUNCTION (_HRESULT_TYPEDEF_(0x87AF0413L))
value SQLITE_E_CONSTRAINT_NOTNULL (_HRESULT_TYPEDEF_(0x87AF0513L))
value SQLITE_E_CONSTRAINT_PRIMARYKEY (_HRESULT_TYPEDEF_(0x87AF0613L))
value SQLITE_E_CONSTRAINT_ROWID (_HRESULT_TYPEDEF_(0x87AF0A13L))
value SQLITE_E_CONSTRAINT_TRIGGER (_HRESULT_TYPEDEF_(0x87AF0713L))
value SQLITE_E_CONSTRAINT_UNIQUE (_HRESULT_TYPEDEF_(0x87AF0813L))
value SQLITE_E_CONSTRAINT_VTAB (_HRESULT_TYPEDEF_(0x87AF0913L))
value SQLITE_E_CORRUPT (_HRESULT_TYPEDEF_(0x87AF000BL))
value SQLITE_E_CORRUPT_VTAB (_HRESULT_TYPEDEF_(0x87AF010BL))
value SQLITE_E_DONE (_HRESULT_TYPEDEF_(0x87AF0065L))
value SQLITE_E_EMPTY (_HRESULT_TYPEDEF_(0x87AF0010L))
value SQLITE_E_ERROR (_HRESULT_TYPEDEF_(0x87AF0001L))
value SQLITE_E_FORMAT (_HRESULT_TYPEDEF_(0x87AF0018L))
value SQLITE_E_FULL (_HRESULT_TYPEDEF_(0x87AF000DL))
value SQLITE_E_INTERNAL (_HRESULT_TYPEDEF_(0x87AF0002L))
value SQLITE_E_INTERRUPT (_HRESULT_TYPEDEF_(0x87AF0009L))
value SQLITE_E_IOERR (_HRESULT_TYPEDEF_(0x87AF000AL))
value SQLITE_E_IOERR_ACCESS (_HRESULT_TYPEDEF_(0x87AF0D0AL))
value SQLITE_E_IOERR_AUTH (_HRESULT_TYPEDEF_(0x87AF1A03L))
value SQLITE_E_IOERR_BLOCKED (_HRESULT_TYPEDEF_(0x87AF0B0AL))
value SQLITE_E_IOERR_CHECKRESERVEDLOCK (_HRESULT_TYPEDEF_(0x87AF0E0AL))
value SQLITE_E_IOERR_CLOSE (_HRESULT_TYPEDEF_(0x87AF100AL))
value SQLITE_E_IOERR_CONVPATH (_HRESULT_TYPEDEF_(0x87AF1A0AL))
value SQLITE_E_IOERR_DELETE (_HRESULT_TYPEDEF_(0x87AF0A0AL))
value SQLITE_E_IOERR_DELETE_NOENT (_HRESULT_TYPEDEF_(0x87AF170AL))
value SQLITE_E_IOERR_DIR_CLOSE (_HRESULT_TYPEDEF_(0x87AF110AL))
value SQLITE_E_IOERR_DIR_FSYNC (_HRESULT_TYPEDEF_(0x87AF050AL))
value SQLITE_E_IOERR_FSTAT (_HRESULT_TYPEDEF_(0x87AF070AL))
value SQLITE_E_IOERR_FSYNC (_HRESULT_TYPEDEF_(0x87AF040AL))
value SQLITE_E_IOERR_GETTEMPPATH (_HRESULT_TYPEDEF_(0x87AF190AL))
value SQLITE_E_IOERR_LOCK (_HRESULT_TYPEDEF_(0x87AF0F0AL))
value SQLITE_E_IOERR_MMAP (_HRESULT_TYPEDEF_(0x87AF180AL))
value SQLITE_E_IOERR_NOMEM (_HRESULT_TYPEDEF_(0x87AF0C0AL))
value SQLITE_E_IOERR_RDLOCK (_HRESULT_TYPEDEF_(0x87AF090AL))
value SQLITE_E_IOERR_READ (_HRESULT_TYPEDEF_(0x87AF010AL))
value SQLITE_E_IOERR_SEEK (_HRESULT_TYPEDEF_(0x87AF160AL))
value SQLITE_E_IOERR_SHMLOCK (_HRESULT_TYPEDEF_(0x87AF140AL))
value SQLITE_E_IOERR_SHMMAP (_HRESULT_TYPEDEF_(0x87AF150AL))
value SQLITE_E_IOERR_SHMOPEN (_HRESULT_TYPEDEF_(0x87AF120AL))
value SQLITE_E_IOERR_SHMSIZE (_HRESULT_TYPEDEF_(0x87AF130AL))
value SQLITE_E_IOERR_SHORT_READ (_HRESULT_TYPEDEF_(0x87AF020AL))
value SQLITE_E_IOERR_TRUNCATE (_HRESULT_TYPEDEF_(0x87AF060AL))
value SQLITE_E_IOERR_UNLOCK (_HRESULT_TYPEDEF_(0x87AF080AL))
value SQLITE_E_IOERR_VNODE (_HRESULT_TYPEDEF_(0x87AF1A02L))
value SQLITE_E_IOERR_WRITE (_HRESULT_TYPEDEF_(0x87AF030AL))
value SQLITE_E_LOCKED (_HRESULT_TYPEDEF_(0x87AF0006L))
value SQLITE_E_LOCKED_SHAREDCACHE (_HRESULT_TYPEDEF_(0x87AF0106L))
value SQLITE_E_MISMATCH (_HRESULT_TYPEDEF_(0x87AF0014L))
value SQLITE_E_MISUSE (_HRESULT_TYPEDEF_(0x87AF0015L))
value SQLITE_E_NOLFS (_HRESULT_TYPEDEF_(0x87AF0016L))
value SQLITE_E_NOMEM (_HRESULT_TYPEDEF_(0x87AF0007L))
value SQLITE_E_NOTADB (_HRESULT_TYPEDEF_(0x87AF001AL))
value SQLITE_E_NOTFOUND (_HRESULT_TYPEDEF_(0x87AF000CL))
value SQLITE_E_NOTICE (_HRESULT_TYPEDEF_(0x87AF001BL))
value SQLITE_E_NOTICE_RECOVER_ROLLBACK (_HRESULT_TYPEDEF_(0x87AF021BL))
value SQLITE_E_NOTICE_RECOVER_WAL (_HRESULT_TYPEDEF_(0x87AF011BL))
value SQLITE_E_PERM (_HRESULT_TYPEDEF_(0x87AF0003L))
value SQLITE_E_PROTOCOL (_HRESULT_TYPEDEF_(0x87AF000FL))
value SQLITE_E_RANGE (_HRESULT_TYPEDEF_(0x87AF0019L))
value SQLITE_E_READONLY (_HRESULT_TYPEDEF_(0x87AF0008L))
value SQLITE_E_READONLY_CANTLOCK (_HRESULT_TYPEDEF_(0x87AF0208L))
value SQLITE_E_READONLY_DBMOVED (_HRESULT_TYPEDEF_(0x87AF0408L))
value SQLITE_E_READONLY_RECOVERY (_HRESULT_TYPEDEF_(0x87AF0108L))
value SQLITE_E_READONLY_ROLLBACK (_HRESULT_TYPEDEF_(0x87AF0308L))
value SQLITE_E_ROW (_HRESULT_TYPEDEF_(0x87AF0064L))
value SQLITE_E_SCHEMA (_HRESULT_TYPEDEF_(0x87AF0011L))
value SQLITE_E_TOOBIG (_HRESULT_TYPEDEF_(0x87AF0012L))
value SQLITE_E_WARNING (_HRESULT_TYPEDEF_(0x87AF001CL))
value SQLITE_E_WARNING_AUTOINDEX (_HRESULT_TYPEDEF_(0x87AF011CL))
value SRB_TYPE_SCSI_REQUEST_BLOCK (0)
value SRB_TYPE_STORAGE_REQUEST_BLOCK (1)
value SRCAND ((DWORD)0x008800C6)
value SRCCOPY ((DWORD)0x00CC0020)
value SRCERASE ((DWORD)0x00440328)
value SRCINVERT ((DWORD)0x00660046)
value SRCPAINT ((DWORD)0x00EE0086)
value SRWLOCK_INIT (RTL_SRWLOCK_INIT)
value SSF_AVAILABLE (0x00000002)
value SSF_INDICATOR (0x00000004)
value SSF_SOUNDSENTRYON (0x00000001)
value SSGF_DISPLAY (3)
value SSGF_NONE (0)
value SSL_HPKP_HEADER_COUNT (2)
value SSL_HPKP_PKP_HEADER_INDEX (0)
value SSL_HPKP_PKP_RO_HEADER_INDEX (1)
value SSL_KEY_PIN_ERROR_TEXT_LENGTH (512)
value SSTF_BORDER (2)
value SSTF_CHARS (1)
value SSTF_DISPLAY (3)
value SSTF_NONE (0)
value SSWF_CUSTOM (4)
value SSWF_DISPLAY (3)
value SSWF_NONE (0)
value SSWF_TITLE (1)
value SSWF_WINDOW (2)
value SS_BITMAP (0x0000000EL)
value SS_BLACKFRAME (0x00000007L)
value SS_BLACKRECT (0x00000004L)
value SS_CENTER (0x00000001L)
value SS_CENTERIMAGE (0x00000200L)
value SS_EDITCONTROL (0x00002000L)
value SS_ELLIPSISMASK (0x0000C000L)
value SS_ENDELLIPSIS (0x00004000L)
value SS_ENHMETAFILE (0x0000000FL)
value SS_ETCHEDFRAME (0x00000012L)
value SS_ETCHEDHORZ (0x00000010L)
value SS_ETCHEDVERT (0x00000011L)
value SS_GRAYFRAME (0x00000008L)
value SS_GRAYRECT (0x00000005L)
value SS_ICON (0x00000003L)
value SS_LEFT (0x00000000L)
value SS_LEFTNOWORDWRAP (0x0000000CL)
value SS_NOPREFIX (0x00000080L)
value SS_NOTIFY (0x00000100L)
value SS_OWNERDRAW (0x0000000DL)
value SS_PATHELLIPSIS (0x00008000L)
value SS_REALSIZECONTROL (0x00000040L)
value SS_REALSIZEIMAGE (0x00000800L)
value SS_RIGHT (0x00000002L)
value SS_RIGHTJUST (0x00000400L)
value SS_SIMPLE (0x0000000BL)
value SS_SUNKEN (0x00001000L)
value SS_TYPEMASK (0x0000001FL)
value SS_USERITEM (0x0000000AL)
value SS_WHITEFRAME (0x00000009L)
value SS_WHITERECT (0x00000006L)
value SS_WORDELLIPSIS (0x0000C000L)
value STACK_SIZE_PARAM_IS_A_RESERVATION (0x00010000)
value STANDARD_RIGHTS_ALL ((0x001F0000L))
value STANDARD_RIGHTS_EXECUTE ((READ_CONTROL))
value STANDARD_RIGHTS_READ ((READ_CONTROL))
value STANDARD_RIGHTS_REQUIRED ((0x000F0000L))
value STANDARD_RIGHTS_WRITE ((READ_CONTROL))
value STARTDOC (10)
value STARTF_FORCEOFFFEEDBACK (0x00000080)
value STARTF_FORCEONFEEDBACK (0x00000040)
value STARTF_HOLOGRAPHIC (0x00040000)
value STARTF_PREVENTPINNING (0x00002000)
value STARTF_RUNFULLSCREEN (0x00000020)
value STARTF_TITLEISAPPID (0x00001000)
value STARTF_TITLEISLINKNAME (0x00000800)
value STARTF_UNTRUSTEDSOURCE (0x00008000)
value STARTF_USECOUNTCHARS (0x00000008)
value STARTF_USEFILLATTRIBUTE (0x00000010)
value STARTF_USEHOTKEY (0x00000200)
value STARTF_USEPOSITION (0x00000004)
value STARTF_USESHOWWINDOW (0x00000001)
value STARTF_USESIZE (0x00000002)
value STARTF_USESTDHANDLES (0x00000100)
value START_PAGE_GENERAL (0xffffffff)
value STATEREPOSITORY_ERROR_CACHE_CORRUPTED (_HRESULT_TYPEDEF_(0x80670012L))
value STATEREPOSITORY_ERROR_DICTIONARY_CORRUPTED (_HRESULT_TYPEDEF_(0x80670005L))
value STATEREPOSITORY_E_BLOCKED (_HRESULT_TYPEDEF_(0x80670006L))
value STATEREPOSITORY_E_BUSY_RECOVERY_RETRY (_HRESULT_TYPEDEF_(0x80670008L))
value STATEREPOSITORY_E_BUSY_RECOVERY_TIMEOUT_EXCEEDED (_HRESULT_TYPEDEF_(0x8067000DL))
value STATEREPOSITORY_E_BUSY_RETRY (_HRESULT_TYPEDEF_(0x80670007L))
value STATEREPOSITORY_E_BUSY_TIMEOUT_EXCEEDED (_HRESULT_TYPEDEF_(0x8067000CL))
value STATEREPOSITORY_E_CACHE_NOT_INIITALIZED (_HRESULT_TYPEDEF_(0x80670015L))
value STATEREPOSITORY_E_CONCURRENCY_LOCKING_FAILURE (_HRESULT_TYPEDEF_(0x80670001L))
value STATEREPOSITORY_E_CONFIGURATION_INVALID (_HRESULT_TYPEDEF_(0x80670003L))
value STATEREPOSITORY_E_DEPENDENCY_NOT_RESOLVED (_HRESULT_TYPEDEF_(0x80670016L))
value STATEREPOSITORY_E_LOCKED_RETRY (_HRESULT_TYPEDEF_(0x80670009L))
value STATEREPOSITORY_E_LOCKED_SHAREDCACHE_RETRY (_HRESULT_TYPEDEF_(0x8067000AL))
value STATEREPOSITORY_E_LOCKED_SHAREDCACHE_TIMEOUT_EXCEEDED (_HRESULT_TYPEDEF_(0x8067000FL))
value STATEREPOSITORY_E_LOCKED_TIMEOUT_EXCEEDED (_HRESULT_TYPEDEF_(0x8067000EL))
value STATEREPOSITORY_E_SERVICE_STOP_IN_PROGRESS (_HRESULT_TYPEDEF_(0x80670010L))
value STATEREPOSITORY_E_STATEMENT_INPROGRESS (_HRESULT_TYPEDEF_(0x80670002L))
value STATEREPOSITORY_E_TRANSACTION_REQUIRED (_HRESULT_TYPEDEF_(0x8067000BL))
value STATEREPOSITORY_E_UNKNOWN_SCHEMA_VERSION (_HRESULT_TYPEDEF_(0x80670004L))
value STATEREPOSITORY_TRANSACTION_CALLER_ID_CHANGED (_HRESULT_TYPEDEF_(0x00670013L))
value STATEREPOSITORY_TRANSACTION_IN_PROGRESS (_HRESULT_TYPEDEF_(0x80670014L))
value STATEREPOSTORY_E_NESTED_TRANSACTION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80670011L))
value STATE_SYSTEM_ALERT_HIGH (0x10000000)
value STATE_SYSTEM_ALERT_LOW (0x04000000)
value STATE_SYSTEM_ALERT_MEDIUM (0x08000000)
value STATE_SYSTEM_ANIMATED (0x00004000)
value STATE_SYSTEM_BUSY (0x00000800)
value STATE_SYSTEM_CHECKED (0x00000010)
value STATE_SYSTEM_COLLAPSED (0x00000400)
value STATE_SYSTEM_DEFAULT (0x00000100)
value STATE_SYSTEM_EXPANDED (0x00000200)
value STATE_SYSTEM_EXTSELECTABLE (0x02000000)
value STATE_SYSTEM_FLOATING (0x00001000)
value STATE_SYSTEM_FOCUSABLE (0x00100000)
value STATE_SYSTEM_FOCUSED (0x00000004)
value STATE_SYSTEM_HOTTRACKED (0x00000080)
value STATE_SYSTEM_INDETERMINATE (STATE_SYSTEM_MIXED)
value STATE_SYSTEM_INVISIBLE (0x00008000)
value STATE_SYSTEM_LINKED (0x00400000)
value STATE_SYSTEM_MARQUEED (0x00002000)
value STATE_SYSTEM_MIXED (0x00000020)
value STATE_SYSTEM_MOVEABLE (0x00040000)
value STATE_SYSTEM_MULTISELECTABLE (0x01000000)
value STATE_SYSTEM_OFFSCREEN (0x00010000)
value STATE_SYSTEM_PRESSED (0x00000008)
value STATE_SYSTEM_PROTECTED (0x20000000)
value STATE_SYSTEM_READONLY (0x00000040)
value STATE_SYSTEM_SELECTABLE (0x00200000)
value STATE_SYSTEM_SELECTED (0x00000002)
value STATE_SYSTEM_SELFVOICING (0x00080000)
value STATE_SYSTEM_SIZEABLE (0x00020000)
value STATE_SYSTEM_TRAVERSED (0x00800000)
value STATE_SYSTEM_UNAVAILABLE (0x00000001)
value STATE_SYSTEM_VALID (0x3FFFFFFF)
value STATUS_ACCESS_VIOLATION (((DWORD )0xC0000005L))
value STATUS_ALREADY_REGISTERED (((DWORD )0xC0000718L))
value STATUS_ARRAY_BOUNDS_EXCEEDED (((DWORD )0xC000008CL))
value STATUS_ASSERTION_FAILURE (((DWORD )0xC0000420L))
value STATUS_BREAKPOINT (((DWORD )0x80000003L))
value STATUS_CONTROL_C_EXIT (((DWORD )0xC000013AL))
value STATUS_CONTROL_STACK_VIOLATION (((DWORD )0xC00001B2L))
value STATUS_DATATYPE_MISALIGNMENT (((DWORD )0x80000002L))
value STATUS_DLL_INIT_FAILED (((DWORD )0xC0000142L))
value STATUS_DLL_NOT_FOUND (((DWORD )0xC0000135L))
value STATUS_ENCLAVE_VIOLATION (((DWORD )0xC00004A2L))
value STATUS_ENTRYPOINT_NOT_FOUND (((DWORD )0xC0000139L))
value STATUS_FATAL_APP_EXIT (((DWORD )0x40000015L))
value STATUS_FLOAT_DENORMAL_OPERAND (((DWORD )0xC000008DL))
value STATUS_FLOAT_DIVIDE_BY_ZERO (((DWORD )0xC000008EL))
value STATUS_FLOAT_INEXACT_RESULT (((DWORD )0xC000008FL))
value STATUS_FLOAT_INVALID_OPERATION (((DWORD )0xC0000090L))
value STATUS_FLOAT_MULTIPLE_FAULTS (((DWORD )0xC00002B4L))
value STATUS_FLOAT_MULTIPLE_TRAPS (((DWORD )0xC00002B5L))
value STATUS_FLOAT_OVERFLOW (((DWORD )0xC0000091L))
value STATUS_FLOAT_STACK_CHECK (((DWORD )0xC0000092L))
value STATUS_FLOAT_UNDERFLOW (((DWORD )0xC0000093L))
value STATUS_GUARD_PAGE_VIOLATION (((DWORD )0x80000001L))
value STATUS_HEAP_CORRUPTION (((DWORD )0xC0000374L))
value STATUS_ILLEGAL_INSTRUCTION (((DWORD )0xC000001DL))
value STATUS_INTEGER_DIVIDE_BY_ZERO (((DWORD )0xC0000094L))
value STATUS_INTEGER_OVERFLOW (((DWORD )0xC0000095L))
value STATUS_INTERRUPTED (((DWORD )0xC0000515L))
value STATUS_INVALID_CRUNTIME_PARAMETER (((DWORD )0xC0000417L))
value STATUS_INVALID_DISPOSITION (((DWORD )0xC0000026L))
value STATUS_INVALID_HANDLE (((DWORD )0xC0000008L))
value STATUS_INVALID_PARAMETER (((DWORD )0xC000000DL))
value STATUS_IN_PAGE_ERROR (((DWORD )0xC0000006L))
value STATUS_LONGJUMP (((DWORD )0x80000026L))
value STATUS_NONCONTINUABLE_EXCEPTION (((DWORD )0xC0000025L))
value STATUS_NO_MEMORY (((DWORD )0xC0000017L))
value STATUS_ORDINAL_NOT_FOUND (((DWORD )0xC0000138L))
value STATUS_PENDING (((DWORD )0x00000103L))
value STATUS_PRIVILEGED_INSTRUCTION (((DWORD )0xC0000096L))
value STATUS_REG_NAT_CONSUMPTION (((DWORD )0xC00002C9L))
value STATUS_SEGMENT_NOTIFICATION (((DWORD )0x40000005L))
value STATUS_SINGLE_STEP (((DWORD )0x80000004L))
value STATUS_STACK_BUFFER_OVERRUN (((DWORD )0xC0000409L))
value STATUS_STACK_OVERFLOW (((DWORD )0xC00000FDL))
value STATUS_SXS_EARLY_DEACTIVATION (((DWORD )0xC015000FL))
value STATUS_SXS_INVALID_DEACTIVATION (((DWORD )0xC0150010L))
value STATUS_THREAD_NOT_RUNNING (((DWORD )0xC0000516L))
value STATUS_TIMEOUT (((DWORD )0x00000102L))
value STATUS_UNWIND_CONSOLIDATE (((DWORD )0x80000029L))
value STATUS_USER_APC (((DWORD )0x000000C0L))
value STDAPI (EXTERN_C HRESULT STDAPICALLTYPE)
value STDAPIV (EXTERN_C HRESULT STDAPIVCALLTYPE)
value STDMETHODIMP (HRESULT STDMETHODCALLTYPE)
value STDMETHODIMPV (HRESULT STDMETHODVCALLTYPE)
value STDOLE_LCID (0x0000)
value STDOLE_MAJORVERNUM (0x1)
value STDOLE_MINORVERNUM (0x0)
value STD_ERROR_HANDLE (((DWORD)-12))
value STD_INPUT_HANDLE (((DWORD)-10))
value STD_OUTPUT_HANDLE (((DWORD)-11))
value STGFMT_ANY (4)
value STGFMT_DOCFILE (5)
value STGFMT_DOCUMENT (0)
value STGFMT_FILE (3)
value STGFMT_NATIVE (1)
value STGFMT_STORAGE (0)
value STGM_CONVERT (0x00020000L)
value STGM_CREATE (0x00001000L)
value STGM_DELETEONRELEASE (0x04000000L)
value STGM_DIRECT (0x00000000L)
value STGM_DIRECT_SWMR (0x00400000L)
value STGM_FAILIFTHERE (0x00000000L)
value STGM_NOSCRATCH (0x00100000L)
value STGM_NOSNAPSHOT (0x00200000L)
value STGM_PRIORITY (0x00040000L)
value STGM_READ (0x00000000L)
value STGM_READWRITE (0x00000002L)
value STGM_SHARE_DENY_NONE (0x00000040L)
value STGM_SHARE_DENY_READ (0x00000030L)
value STGM_SHARE_DENY_WRITE (0x00000020L)
value STGM_SHARE_EXCLUSIVE (0x00000010L)
value STGM_SIMPLE (0x08000000L)
value STGM_TRANSACTED (0x00010000L)
value STGM_WRITE (0x00000001L)
value STGOPTIONS_VERSION (2)
value STGTY_REPEAT (0x00000100L)
value STG_E_ABNORMALAPIEXIT (_HRESULT_TYPEDEF_(0x800300FAL))
value STG_E_ACCESSDENIED (_HRESULT_TYPEDEF_(0x80030005L))
value STG_E_BADBASEADDRESS (_HRESULT_TYPEDEF_(0x80030110L))
value STG_E_CANTSAVE (_HRESULT_TYPEDEF_(0x80030103L))
value STG_E_CSS_AUTHENTICATION_FAILURE (_HRESULT_TYPEDEF_(0x80030306L))
value STG_E_CSS_KEY_NOT_ESTABLISHED (_HRESULT_TYPEDEF_(0x80030308L))
value STG_E_CSS_KEY_NOT_PRESENT (_HRESULT_TYPEDEF_(0x80030307L))
value STG_E_CSS_REGION_MISMATCH (_HRESULT_TYPEDEF_(0x8003030AL))
value STG_E_CSS_SCRAMBLED_SECTOR (_HRESULT_TYPEDEF_(0x80030309L))
value STG_E_DEVICE_UNRESPONSIVE (_HRESULT_TYPEDEF_(0x8003020AL))
value STG_E_DISKISWRITEPROTECTED (_HRESULT_TYPEDEF_(0x80030013L))
value STG_E_DOCFILECORRUPT (_HRESULT_TYPEDEF_(0x80030109L))
value STG_E_DOCFILETOOLARGE (_HRESULT_TYPEDEF_(0x80030111L))
value STG_E_EXTANTMARSHALLINGS (_HRESULT_TYPEDEF_(0x80030108L))
value STG_E_FILEALREADYEXISTS (_HRESULT_TYPEDEF_(0x80030050L))
value STG_E_FILENOTFOUND (_HRESULT_TYPEDEF_(0x80030002L))
value STG_E_FIRMWARE_IMAGE_INVALID (_HRESULT_TYPEDEF_(0x80030209L))
value STG_E_FIRMWARE_SLOT_INVALID (_HRESULT_TYPEDEF_(0x80030208L))
value STG_E_INCOMPLETE (_HRESULT_TYPEDEF_(0x80030201L))
value STG_E_INSUFFICIENTMEMORY (_HRESULT_TYPEDEF_(0x80030008L))
value STG_E_INUSE (_HRESULT_TYPEDEF_(0x80030100L))
value STG_E_INVALIDFLAG (_HRESULT_TYPEDEF_(0x800300FFL))
value STG_E_INVALIDFUNCTION (_HRESULT_TYPEDEF_(0x80030001L))
value STG_E_INVALIDHANDLE (_HRESULT_TYPEDEF_(0x80030006L))
value STG_E_INVALIDHEADER (_HRESULT_TYPEDEF_(0x800300FBL))
value STG_E_INVALIDNAME (_HRESULT_TYPEDEF_(0x800300FCL))
value STG_E_INVALIDPARAMETER (_HRESULT_TYPEDEF_(0x80030057L))
value STG_E_INVALIDPOINTER (_HRESULT_TYPEDEF_(0x80030009L))
value STG_E_LOCKVIOLATION (_HRESULT_TYPEDEF_(0x80030021L))
value STG_E_MEDIUMFULL (_HRESULT_TYPEDEF_(0x80030070L))
value STG_E_NOMOREFILES (_HRESULT_TYPEDEF_(0x80030012L))
value STG_E_NOTCURRENT (_HRESULT_TYPEDEF_(0x80030101L))
value STG_E_NOTFILEBASEDSTORAGE (_HRESULT_TYPEDEF_(0x80030107L))
value STG_E_NOTSIMPLEFORMAT (_HRESULT_TYPEDEF_(0x80030112L))
value STG_E_OLDDLL (_HRESULT_TYPEDEF_(0x80030105L))
value STG_E_OLDFORMAT (_HRESULT_TYPEDEF_(0x80030104L))
value STG_E_PATHNOTFOUND (_HRESULT_TYPEDEF_(0x80030003L))
value STG_E_PROPSETMISMATCHED (_HRESULT_TYPEDEF_(0x800300F0L))
value STG_E_READFAULT (_HRESULT_TYPEDEF_(0x8003001EL))
value STG_E_RESETS_EXHAUSTED (_HRESULT_TYPEDEF_(0x8003030BL))
value STG_E_REVERTED (_HRESULT_TYPEDEF_(0x80030102L))
value STG_E_SEEKERROR (_HRESULT_TYPEDEF_(0x80030019L))
value STG_E_SHAREREQUIRED (_HRESULT_TYPEDEF_(0x80030106L))
value STG_E_SHAREVIOLATION (_HRESULT_TYPEDEF_(0x80030020L))
value STG_E_STATUS_COPY_PROTECTION_FAILURE (_HRESULT_TYPEDEF_(0x80030305L))
value STG_E_TERMINATED (_HRESULT_TYPEDEF_(0x80030202L))
value STG_E_TOOMANYOPENFILES (_HRESULT_TYPEDEF_(0x80030004L))
value STG_E_UNIMPLEMENTEDFUNCTION (_HRESULT_TYPEDEF_(0x800300FEL))
value STG_E_UNKNOWN (_HRESULT_TYPEDEF_(0x800300FDL))
value STG_E_WRITEFAULT (_HRESULT_TYPEDEF_(0x8003001DL))
value STG_LAYOUT_INTERLEAVED (0x00000001L)
value STG_LAYOUT_SEQUENTIAL (0x00000000L)
value STG_S_BLOCK (_HRESULT_TYPEDEF_(0x00030201L))
value STG_S_CANNOTCONSOLIDATE (_HRESULT_TYPEDEF_(0x00030206L))
value STG_S_CONSOLIDATIONFAILED (_HRESULT_TYPEDEF_(0x00030205L))
value STG_S_CONVERTED (_HRESULT_TYPEDEF_(0x00030200L))
value STG_S_MONITORING (_HRESULT_TYPEDEF_(0x00030203L))
value STG_S_MULTIPLEOPENS (_HRESULT_TYPEDEF_(0x00030204L))
value STG_S_POWER_CYCLE_REQUIRED (_HRESULT_TYPEDEF_(0x00030207L))
value STG_S_RETRYNOW (_HRESULT_TYPEDEF_(0x00030202L))
value STG_TOEND (0xFFFFFFFFL)
value STILL_ACTIVE (STATUS_PENDING)
value STKFORCEINLINE (FORCEINLINE)
value STM_GETICON (0x0171)
value STM_GETIMAGE (0x0173)
value STM_MSGMAX (0x0174)
value STM_SETICON (0x0170)
value STM_SETIMAGE (0x0172)
value STN_CLICKED (0)
value STN_DBLCLK (1)
value STN_DISABLE (3)
value STN_ENABLE (2)
value STOCK_LAST (19)
value STORAGE_ATTRIBUTE_ASYNC_EVENT_NOTIFICATION (0x10)
value STORAGE_ATTRIBUTE_BLOCK_IO (0x02)
value STORAGE_ATTRIBUTE_BYTE_ADDRESSABLE_IO (0x01)
value STORAGE_ATTRIBUTE_DYNAMIC_PERSISTENCE (0x04)
value STORAGE_ATTRIBUTE_PERF_SIZE_INDEPENDENT (0x20)
value STORAGE_ATTRIBUTE_VOLATILE (0x08)
value STORAGE_COMPONENT_ROLE_CACHE (0x00000001)
value STORAGE_COMPONENT_ROLE_DATA (0x00000004)
value STORAGE_COMPONENT_ROLE_TIERING (0x00000002)
value STORAGE_DEVICE_FLAGS_RANDOM_DEVICEGUID_REASON_CONFLICT (0x1)
value STORAGE_DEVICE_FLAGS_RANDOM_DEVICEGUID_REASON_NOHWID (0x2)
value STORAGE_DEVICE_MAX_OPERATIONAL_STATUS (16)
value STORAGE_DEVICE_NUMA_NODE_UNKNOWN (MAXDWORD)
value STORAGE_DIAGNOSTIC_FLAG_ADAPTER_REQUEST (0x00000001)
value STORAGE_EVENT_ALL ((STORAGE_EVENT_MEDIA_STATUS | STORAGE_EVENT_DEVICE_STATUS | STORAGE_EVENT_DEVICE_OPERATION))
value STORAGE_EVENT_DEVICE_OPERATION (0x0000000000000004)
value STORAGE_EVENT_DEVICE_STATUS (0x0000000000000002)
value STORAGE_EVENT_MEDIA_STATUS (0x0000000000000001)
value STORAGE_HW_FIRMWARE_INVALID_SLOT (0xFF)
value STORAGE_HW_FIRMWARE_REQUEST_FLAG_CONTROLLER (0x00000001)
value STORAGE_HW_FIRMWARE_REQUEST_FLAG_FIRST_SEGMENT (0x00000004)
value STORAGE_HW_FIRMWARE_REQUEST_FLAG_LAST_SEGMENT (0x00000002)
value STORAGE_HW_FIRMWARE_REQUEST_FLAG_REPLACE_EXISTING_IMAGE (0x40000000)
value STORAGE_HW_FIRMWARE_REQUEST_FLAG_SWITCH_TO_EXISTING_FIRMWARE (0x80000000)
value STORAGE_HW_FIRMWARE_REVISION_LENGTH (16)
value STORAGE_INFO_FLAGS_ALIGNED_DEVICE (0x00000001)
value STORAGE_INFO_FLAGS_PARTITION_ALIGNED_ON_DEVICE (0x00000002)
value STORAGE_OFFLOAD_MAX_TOKEN_LENGTH (512)
value STORAGE_OFFLOAD_READ_RANGE_TRUNCATED (0x00000001)
value STORAGE_OFFLOAD_TOKEN_ID_LENGTH (0x1F8)
value STORAGE_OFFLOAD_TOKEN_INVALID (0x0002)
value STORAGE_OFFLOAD_TOKEN_TYPE_ZERO_DATA (0xFFFF0001)
value STORAGE_OFFLOAD_WRITE_RANGE_TRUNCATED (0x0001)
value STORAGE_PRIORITY_HINT_SUPPORTED (0x0001)
value STORAGE_PROTOCOL_COMMAND_FLAG_ADAPTER_REQUEST (0x80000000)
value STORAGE_PROTOCOL_COMMAND_LENGTH_NVME (0x40)
value STORAGE_PROTOCOL_SPECIFIC_NVME_ADMIN_COMMAND (0x01)
value STORAGE_PROTOCOL_SPECIFIC_NVME_NVM_COMMAND (0x02)
value STORAGE_PROTOCOL_STATUS_BUSY (0x5)
value STORAGE_PROTOCOL_STATUS_DATA_OVERRUN (0x6)
value STORAGE_PROTOCOL_STATUS_ERROR (0x2)
value STORAGE_PROTOCOL_STATUS_INSUFFICIENT_RESOURCES (0x7)
value STORAGE_PROTOCOL_STATUS_INVALID_REQUEST (0x3)
value STORAGE_PROTOCOL_STATUS_NOT_SUPPORTED (0xFF)
value STORAGE_PROTOCOL_STATUS_NO_DEVICE (0x4)
value STORAGE_PROTOCOL_STATUS_PENDING (0x0)
value STORAGE_PROTOCOL_STATUS_SUCCESS (0x1)
value STORAGE_PROTOCOL_STATUS_THROTTLED_REQUEST (0x8)
value STORAGE_PROTOCOL_STRUCTURE_VERSION (0x1)
value STORAGE_RPMB_MINIMUM_RELIABLE_WRITE_SIZE (512)
value STORAGE_TEMPERATURE_THRESHOLD_FLAG_ADAPTER_REQUEST (0x0001)
value STORAGE_TEMPERATURE_VALUE_NOT_REPORTED (0x8000)
value STORAGE_TIER_DESCRIPTION_LENGTH ((512))
value STORAGE_TIER_FLAG_NO_SEEK_PENALTY ((0x00020000))
value STORAGE_TIER_FLAG_PARITY ((0x00800000))
value STORAGE_TIER_FLAG_READ_CACHE ((0x00400000))
value STORAGE_TIER_FLAG_SMR ((0x01000000))
value STORAGE_TIER_FLAG_WRITE_BACK_CACHE ((0x00200000))
value STORAGE_TIER_NAME_LENGTH ((256))
value STORATTRIBUTE_MANAGEMENT_STATE (1)
value STORATTRIBUTE_NONE (0)
value STORE_ERROR_LICENSE_REVOKED (15864)
value STORE_ERROR_PENDING_COM_TRANSACTION (15863)
value STORE_ERROR_UNLICENSED (15861)
value STORE_ERROR_UNLICENSED_USER (15862)
value STREAMS_ASSOCIATE_ID_CLEAR ((0x1))
value STREAMS_ASSOCIATE_ID_SET ((0x2))
value STREAMS_INVALID_ID ((0))
value STREAMS_MAX_ID ((MAXWORD ))
value STREAM_CLEAR_ENCRYPTION (0x00000004)
value STREAM_CONTAINS_GHOSTED_FILE_EXTENTS (0x00000010)
value STREAM_CONTAINS_PROPERTIES (0x00000004)
value STREAM_CONTAINS_SECURITY (0x00000002)
value STREAM_EXTENT_ENTRY_ALL_EXTENTS ((0x00000002))
value STREAM_EXTENT_ENTRY_AS_RETRIEVAL_POINTERS ((0x00000001))
value STREAM_LAYOUT_ENTRY_HAS_INFORMATION ((0x00000010))
value STREAM_LAYOUT_ENTRY_IMMOVABLE ((0x00000001))
value STREAM_LAYOUT_ENTRY_NO_CLUSTERS_ALLOCATED ((0x00000008))
value STREAM_LAYOUT_ENTRY_PINNED ((0x00000002))
value STREAM_LAYOUT_ENTRY_RESIDENT ((0x00000004))
value STREAM_MODIFIED_WHEN_READ (0x00000001)
value STREAM_NORMAL_ATTRIBUTE (0x00000000)
value STREAM_SET_ENCRYPTION (0x00000003)
value STREAM_SPARSE_ATTRIBUTE (0x00000008)
value STRETCHBLT (2048)
value STRETCH_ANDSCANS (BLACKONWHITE)
value STRETCH_DELETESCANS (COLORONCOLOR)
value STRETCH_HALFTONE (HALFTONE)
value STRETCH_ORSCANS (WHITEONBLACK)
value STRICT (1)
value STRING_LANGPAIR (0x00000004)
value STRING_MUIDLL (0x00000002)
value STRING_NONE (0x00000001)
value STRUNCATE (80)
value STYLE_DESCRIPTION_SIZE (32)
value ST_ADVISE (0x0002)
value ST_BLOCKED (0x0008)
value ST_BLOCKNEXT (0x0080)
value ST_CLIENT (0x0010)
value ST_CONNECTED (0x0001)
value ST_INLIST (0x0040)
value ST_ISLOCAL (0x0004)
value ST_ISSELF (0x0100)
value ST_TERMINATED (0x0020)
value SUBLANG_AFRIKAANS_SOUTH_AFRICA (0x01)
value SUBLANG_ALBANIAN_ALBANIA (0x01)
value SUBLANG_ALSATIAN_FRANCE (0x01)
value SUBLANG_AMHARIC_ETHIOPIA (0x01)
value SUBLANG_ARABIC_ALGERIA (0x05)
value SUBLANG_ARABIC_BAHRAIN (0x0f)
value SUBLANG_ARABIC_EGYPT (0x03)
value SUBLANG_ARABIC_IRAQ (0x02)
value SUBLANG_ARABIC_JORDAN (0x0b)
value SUBLANG_ARABIC_KUWAIT (0x0d)
value SUBLANG_ARABIC_LEBANON (0x0c)
value SUBLANG_ARABIC_LIBYA (0x04)
value SUBLANG_ARABIC_MOROCCO (0x06)
value SUBLANG_ARABIC_OMAN (0x08)
value SUBLANG_ARABIC_QATAR (0x10)
value SUBLANG_ARABIC_SAUDI_ARABIA (0x01)
value SUBLANG_ARABIC_SYRIA (0x0a)
value SUBLANG_ARABIC_TUNISIA (0x07)
value SUBLANG_ARABIC_UAE (0x0e)
value SUBLANG_ARABIC_YEMEN (0x09)
value SUBLANG_ARMENIAN_ARMENIA (0x01)
value SUBLANG_ASSAMESE_INDIA (0x01)
value SUBLANG_AZERBAIJANI_AZERBAIJAN_CYRILLIC (0x02)
value SUBLANG_AZERBAIJANI_AZERBAIJAN_LATIN (0x01)
value SUBLANG_AZERI_CYRILLIC (0x02)
value SUBLANG_AZERI_LATIN (0x01)
value SUBLANG_BANGLA_BANGLADESH (0x02)
value SUBLANG_BANGLA_INDIA (0x01)
value SUBLANG_BASHKIR_RUSSIA (0x01)
value SUBLANG_BASQUE_BASQUE (0x01)
value SUBLANG_BELARUSIAN_BELARUS (0x01)
value SUBLANG_BENGALI_BANGLADESH (0x02)
value SUBLANG_BENGALI_INDIA (0x01)
value SUBLANG_BOSNIAN_BOSNIA_HERZEGOVINA_CYRILLIC (0x08)
value SUBLANG_BOSNIAN_BOSNIA_HERZEGOVINA_LATIN (0x05)
value SUBLANG_BRETON_FRANCE (0x01)
value SUBLANG_BULGARIAN_BULGARIA (0x01)
value SUBLANG_CATALAN_CATALAN (0x01)
value SUBLANG_CENTRAL_KURDISH_IRAQ (0x01)
value SUBLANG_CHEROKEE_CHEROKEE (0x01)
value SUBLANG_CHINESE_HONGKONG (0x03)
value SUBLANG_CHINESE_MACAU (0x05)
value SUBLANG_CHINESE_SIMPLIFIED (0x02)
value SUBLANG_CHINESE_SINGAPORE (0x04)
value SUBLANG_CHINESE_TRADITIONAL (0x01)
value SUBLANG_CORSICAN_FRANCE (0x01)
value SUBLANG_CROATIAN_BOSNIA_HERZEGOVINA_LATIN (0x04)
value SUBLANG_CROATIAN_CROATIA (0x01)
value SUBLANG_CUSTOM_DEFAULT (0x03)
value SUBLANG_CUSTOM_UNSPECIFIED (0x04)
value SUBLANG_CZECH_CZECH_REPUBLIC (0x01)
value SUBLANG_DANISH_DENMARK (0x01)
value SUBLANG_DARI_AFGHANISTAN (0x01)
value SUBLANG_DEFAULT (0x01)
value SUBLANG_DIVEHI_MALDIVES (0x01)
value SUBLANG_DUTCH (0x01)
value SUBLANG_DUTCH_BELGIAN (0x02)
value SUBLANG_ENGLISH_AUS (0x03)
value SUBLANG_ENGLISH_BELIZE (0x0a)
value SUBLANG_ENGLISH_CAN (0x04)
value SUBLANG_ENGLISH_CARIBBEAN (0x09)
value SUBLANG_ENGLISH_EIRE (0x06)
value SUBLANG_ENGLISH_INDIA (0x10)
value SUBLANG_ENGLISH_JAMAICA (0x08)
value SUBLANG_ENGLISH_MALAYSIA (0x11)
value SUBLANG_ENGLISH_NZ (0x05)
value SUBLANG_ENGLISH_PHILIPPINES (0x0d)
value SUBLANG_ENGLISH_SINGAPORE (0x12)
value SUBLANG_ENGLISH_SOUTH_AFRICA (0x07)
value SUBLANG_ENGLISH_TRINIDAD (0x0b)
value SUBLANG_ENGLISH_UK (0x02)
value SUBLANG_ENGLISH_US (0x01)
value SUBLANG_ENGLISH_ZIMBABWE (0x0c)
value SUBLANG_ESTONIAN_ESTONIA (0x01)
value SUBLANG_FAEROESE_FAROE_ISLANDS (0x01)
value SUBLANG_FILIPINO_PHILIPPINES (0x01)
value SUBLANG_FINNISH_FINLAND (0x01)
value SUBLANG_FRENCH (0x01)
value SUBLANG_FRENCH_BELGIAN (0x02)
value SUBLANG_FRENCH_CANADIAN (0x03)
value SUBLANG_FRENCH_LUXEMBOURG (0x05)
value SUBLANG_FRENCH_MONACO (0x06)
value SUBLANG_FRENCH_SWISS (0x04)
value SUBLANG_FRISIAN_NETHERLANDS (0x01)
value SUBLANG_FULAH_SENEGAL (0x02)
value SUBLANG_GALICIAN_GALICIAN (0x01)
value SUBLANG_GEORGIAN_GEORGIA (0x01)
value SUBLANG_GERMAN (0x01)
value SUBLANG_GERMAN_AUSTRIAN (0x03)
value SUBLANG_GERMAN_LIECHTENSTEIN (0x05)
value SUBLANG_GERMAN_LUXEMBOURG (0x04)
value SUBLANG_GERMAN_SWISS (0x02)
value SUBLANG_GREEK_GREECE (0x01)
value SUBLANG_GREENLANDIC_GREENLAND (0x01)
value SUBLANG_GUJARATI_INDIA (0x01)
value SUBLANG_HAUSA_NIGERIA_LATIN (0x01)
value SUBLANG_HAWAIIAN_US (0x01)
value SUBLANG_HEBREW_ISRAEL (0x01)
value SUBLANG_HINDI_INDIA (0x01)
value SUBLANG_HUNGARIAN_HUNGARY (0x01)
value SUBLANG_ICELANDIC_ICELAND (0x01)
value SUBLANG_IGBO_NIGERIA (0x01)
value SUBLANG_INDONESIAN_INDONESIA (0x01)
value SUBLANG_INUKTITUT_CANADA (0x01)
value SUBLANG_INUKTITUT_CANADA_LATIN (0x02)
value SUBLANG_IRISH_IRELAND (0x02)
value SUBLANG_ITALIAN (0x01)
value SUBLANG_ITALIAN_SWISS (0x02)
value SUBLANG_JAPANESE_JAPAN (0x01)
value SUBLANG_KANNADA_INDIA (0x01)
value SUBLANG_KASHMIRI_INDIA (0x02)
value SUBLANG_KASHMIRI_SASIA (0x02)
value SUBLANG_KAZAK_KAZAKHSTAN (0x01)
value SUBLANG_KHMER_CAMBODIA (0x01)
value SUBLANG_KICHE_GUATEMALA (0x01)
value SUBLANG_KINYARWANDA_RWANDA (0x01)
value SUBLANG_KONKANI_INDIA (0x01)
value SUBLANG_KOREAN (0x01)
value SUBLANG_KYRGYZ_KYRGYZSTAN (0x01)
value SUBLANG_LAO_LAO (0x01)
value SUBLANG_LATVIAN_LATVIA (0x01)
value SUBLANG_LITHUANIAN (0x01)
value SUBLANG_LOWER_SORBIAN_GERMANY (0x02)
value SUBLANG_LUXEMBOURGISH_LUXEMBOURG (0x01)
value SUBLANG_MACEDONIAN_MACEDONIA (0x01)
value SUBLANG_MALAYALAM_INDIA (0x01)
value SUBLANG_MALAY_BRUNEI_DARUSSALAM (0x02)
value SUBLANG_MALAY_MALAYSIA (0x01)
value SUBLANG_MALTESE_MALTA (0x01)
value SUBLANG_MAORI_NEW_ZEALAND (0x01)
value SUBLANG_MAPUDUNGUN_CHILE (0x01)
value SUBLANG_MARATHI_INDIA (0x01)
value SUBLANG_MOHAWK_MOHAWK (0x01)
value SUBLANG_MONGOLIAN_CYRILLIC_MONGOLIA (0x01)
value SUBLANG_MONGOLIAN_PRC (0x02)
value SUBLANG_NEPALI_INDIA (0x02)
value SUBLANG_NEPALI_NEPAL (0x01)
value SUBLANG_NEUTRAL (0x00)
value SUBLANG_NORWEGIAN_BOKMAL (0x01)
value SUBLANG_NORWEGIAN_NYNORSK (0x02)
value SUBLANG_OCCITAN_FRANCE (0x01)
value SUBLANG_ODIA_INDIA (0x01)
value SUBLANG_ORIYA_INDIA (0x01)
value SUBLANG_PASHTO_AFGHANISTAN (0x01)
value SUBLANG_PERSIAN_IRAN (0x01)
value SUBLANG_POLISH_POLAND (0x01)
value SUBLANG_PORTUGUESE (0x02)
value SUBLANG_PORTUGUESE_BRAZILIAN (0x01)
value SUBLANG_PULAR_SENEGAL (0x02)
value SUBLANG_PUNJABI_INDIA (0x01)
value SUBLANG_PUNJABI_PAKISTAN (0x02)
value SUBLANG_QUECHUA_BOLIVIA (0x01)
value SUBLANG_QUECHUA_ECUADOR (0x02)
value SUBLANG_QUECHUA_PERU (0x03)
value SUBLANG_ROMANIAN_ROMANIA (0x01)
value SUBLANG_ROMANSH_SWITZERLAND (0x01)
value SUBLANG_RUSSIAN_RUSSIA (0x01)
value SUBLANG_SAKHA_RUSSIA (0x01)
value SUBLANG_SAMI_INARI_FINLAND (0x09)
value SUBLANG_SAMI_LULE_NORWAY (0x04)
value SUBLANG_SAMI_LULE_SWEDEN (0x05)
value SUBLANG_SAMI_NORTHERN_FINLAND (0x03)
value SUBLANG_SAMI_NORTHERN_NORWAY (0x01)
value SUBLANG_SAMI_NORTHERN_SWEDEN (0x02)
value SUBLANG_SAMI_SKOLT_FINLAND (0x08)
value SUBLANG_SAMI_SOUTHERN_NORWAY (0x06)
value SUBLANG_SAMI_SOUTHERN_SWEDEN (0x07)
value SUBLANG_SANSKRIT_INDIA (0x01)
value SUBLANG_SCOTTISH_GAELIC (0x01)
value SUBLANG_SERBIAN_BOSNIA_HERZEGOVINA_CYRILLIC (0x07)
value SUBLANG_SERBIAN_BOSNIA_HERZEGOVINA_LATIN (0x06)
value SUBLANG_SERBIAN_CROATIA (0x01)
value SUBLANG_SERBIAN_CYRILLIC (0x03)
value SUBLANG_SERBIAN_LATIN (0x02)
value SUBLANG_SERBIAN_MONTENEGRO_CYRILLIC (0x0c)
value SUBLANG_SERBIAN_MONTENEGRO_LATIN (0x0b)
value SUBLANG_SERBIAN_SERBIA_CYRILLIC (0x0a)
value SUBLANG_SERBIAN_SERBIA_LATIN (0x09)
value SUBLANG_SINDHI_AFGHANISTAN (0x02)
value SUBLANG_SINDHI_INDIA (0x01)
value SUBLANG_SINDHI_PAKISTAN (0x02)
value SUBLANG_SINHALESE_SRI_LANKA (0x01)
value SUBLANG_SLOVAK_SLOVAKIA (0x01)
value SUBLANG_SLOVENIAN_SLOVENIA (0x01)
value SUBLANG_SOTHO_NORTHERN_SOUTH_AFRICA (0x01)
value SUBLANG_SPANISH (0x01)
value SUBLANG_SPANISH_ARGENTINA (0x0b)
value SUBLANG_SPANISH_BOLIVIA (0x10)
value SUBLANG_SPANISH_CHILE (0x0d)
value SUBLANG_SPANISH_COLOMBIA (0x09)
value SUBLANG_SPANISH_COSTA_RICA (0x05)
value SUBLANG_SPANISH_DOMINICAN_REPUBLIC (0x07)
value SUBLANG_SPANISH_ECUADOR (0x0c)
value SUBLANG_SPANISH_EL_SALVADOR (0x11)
value SUBLANG_SPANISH_GUATEMALA (0x04)
value SUBLANG_SPANISH_HONDURAS (0x12)
value SUBLANG_SPANISH_MEXICAN (0x02)
value SUBLANG_SPANISH_MODERN (0x03)
value SUBLANG_SPANISH_NICARAGUA (0x13)
value SUBLANG_SPANISH_PANAMA (0x06)
value SUBLANG_SPANISH_PARAGUAY (0x0f)
value SUBLANG_SPANISH_PERU (0x0a)
value SUBLANG_SPANISH_PUERTO_RICO (0x14)
value SUBLANG_SPANISH_URUGUAY (0x0e)
value SUBLANG_SPANISH_US (0x15)
value SUBLANG_SPANISH_VENEZUELA (0x08)
value SUBLANG_SWAHILI_KENYA (0x01)
value SUBLANG_SWEDISH (0x01)
value SUBLANG_SWEDISH_FINLAND (0x02)
value SUBLANG_SYRIAC_SYRIA (0x01)
value SUBLANG_SYS_DEFAULT (0x02)
value SUBLANG_TAJIK_TAJIKISTAN (0x01)
value SUBLANG_TAMAZIGHT_ALGERIA_LATIN (0x02)
value SUBLANG_TAMAZIGHT_MOROCCO_TIFINAGH (0x04)
value SUBLANG_TAMIL_INDIA (0x01)
value SUBLANG_TAMIL_SRI_LANKA (0x02)
value SUBLANG_TATAR_RUSSIA (0x01)
value SUBLANG_TELUGU_INDIA (0x01)
value SUBLANG_THAI_THAILAND (0x01)
value SUBLANG_TIBETAN_PRC (0x01)
value SUBLANG_TIGRIGNA_ERITREA (0x02)
value SUBLANG_TIGRINYA_ERITREA (0x02)
value SUBLANG_TIGRINYA_ETHIOPIA (0x01)
value SUBLANG_TSWANA_BOTSWANA (0x02)
value SUBLANG_TSWANA_SOUTH_AFRICA (0x01)
value SUBLANG_TURKISH_TURKEY (0x01)
value SUBLANG_TURKMEN_TURKMENISTAN (0x01)
value SUBLANG_UIGHUR_PRC (0x01)
value SUBLANG_UI_CUSTOM_DEFAULT (0x05)
value SUBLANG_UKRAINIAN_UKRAINE (0x01)
value SUBLANG_UPPER_SORBIAN_GERMANY (0x01)
value SUBLANG_URDU_INDIA (0x02)
value SUBLANG_URDU_PAKISTAN (0x01)
value SUBLANG_UZBEK_CYRILLIC (0x02)
value SUBLANG_UZBEK_LATIN (0x01)
value SUBLANG_VALENCIAN_VALENCIA (0x02)
value SUBLANG_VIETNAMESE_VIETNAM (0x01)
value SUBLANG_WELSH_UNITED_KINGDOM (0x01)
value SUBLANG_WOLOF_SENEGAL (0x01)
value SUBLANG_XHOSA_SOUTH_AFRICA (0x01)
value SUBLANG_YAKUT_RUSSIA (0x01)
value SUBLANG_YI_PRC (0x01)
value SUBLANG_YORUBA_NIGERIA (0x01)
value SUBLANG_ZULU_SOUTH_AFRICA (0x01)
value SUBVERSION_MASK (0x000000FF)
value SUCCESSFUL_ACCESS_ACE_FLAG ((0x40))
value SUPPORT_LANG_NUMBER (32)
value SWP_ASYNCWINDOWPOS (0x4000)
value SWP_DEFERERASE (0x2000)
value SWP_DRAWFRAME (SWP_FRAMECHANGED)
value SWP_FRAMECHANGED (0x0020)
value SWP_HIDEWINDOW (0x0080)
value SWP_NOACTIVATE (0x0010)
value SWP_NOCOPYBITS (0x0100)
value SWP_NOMOVE (0x0002)
value SWP_NOOWNERZORDER (0x0200)
value SWP_NOREDRAW (0x0008)
value SWP_NOREPOSITION (SWP_NOOWNERZORDER)
value SWP_NOSENDCHANGING (0x0400)
value SWP_NOSIZE (0x0001)
value SWP_NOZORDER (0x0004)
value SWP_SHOWWINDOW (0x0040)
value SW_ERASE (0x0004)
value SW_FORCEMINIMIZE (11)
value SW_HIDE (0)
value SW_INVALIDATE (0x0002)
value SW_MAX (11)
value SW_MAXIMIZE (3)
value SW_MINIMIZE (6)
value SW_NORMAL (1)
value SW_OTHERUNZOOM (4)
value SW_OTHERZOOM (2)
value SW_PARENTCLOSING (1)
value SW_PARENTOPENING (3)
value SW_RESTORE (9)
value SW_SCROLLCHILDREN (0x0001)
value SW_SHOW (5)
value SW_SHOWDEFAULT (10)
value SW_SHOWMAXIMIZED (3)
value SW_SHOWMINIMIZED (2)
value SW_SHOWMINNOACTIVE (7)
value SW_SHOWNA (8)
value SW_SHOWNOACTIVATE (4)
value SW_SHOWNORMAL (1)
value SW_SMOOTHSCROLL (0x0010)
value SYMBOLIC_LINK_FLAG_ALLOW_UNPRIVILEGED_CREATE ((0x2))
value SYMBOLIC_LINK_FLAG_DIRECTORY ((0x1))
value SYMBOL_CHARSET (2)
value SYMBOL_FONTTYPE (0x80000)
value SYMMETRICWRAPKEYBLOB (0xB)
value SYNCHRONIZATION_BARRIER_FLAGS_BLOCK_ONLY (0x02)
value SYNCHRONIZATION_BARRIER_FLAGS_NO_DELETE (0x04)
value SYNCHRONIZATION_BARRIER_FLAGS_SPIN_ONLY (0x01)
value SYNCHRONIZE ((0x00100000L))
value SYSPAL_ERROR (0)
value SYSPAL_NOSTATIC (2)
value SYSPAL_STATIC (1)
value SYSRGN (4)
value SYSTEM_ACCESS_FILTER_ACE_TYPE ((0x15))
value SYSTEM_ACCESS_FILTER_NOCONSTRAINT_MASK (0xffffffff)
value SYSTEM_ACCESS_FILTER_VALID_MASK (0x00ffffff)
value SYSTEM_ALARM_ACE_TYPE ((0x3))
value SYSTEM_ALARM_CALLBACK_ACE_TYPE ((0xE))
value SYSTEM_ALARM_CALLBACK_OBJECT_ACE_TYPE ((0x10))
value SYSTEM_ALARM_OBJECT_ACE_TYPE ((0x8))
value SYSTEM_AUDIT_ACE_TYPE ((0x2))
value SYSTEM_AUDIT_CALLBACK_ACE_TYPE ((0xD))
value SYSTEM_AUDIT_CALLBACK_OBJECT_ACE_TYPE ((0xF))
value SYSTEM_AUDIT_OBJECT_ACE_TYPE ((0x7))
value SYSTEM_CACHE_ALIGNMENT_SIZE (X86_CACHE_ALIGNMENT_SIZE)
value SYSTEM_CPU_SET_INFORMATION_ALLOCATED (0x2)
value SYSTEM_CPU_SET_INFORMATION_ALLOCATED_TO_TARGET_PROCESS (0x4)
value SYSTEM_CPU_SET_INFORMATION_PARKED (0x1)
value SYSTEM_CPU_SET_INFORMATION_REALTIME (0x8)
value SYSTEM_FIXED_FONT (16)
value SYSTEM_FONT (13)
value SYSTEM_MANDATORY_LABEL_ACE_TYPE ((0x11))
value SYSTEM_MANDATORY_LABEL_NO_EXECUTE_UP (0x4)
value SYSTEM_MANDATORY_LABEL_NO_READ_UP (0x2)
value SYSTEM_MANDATORY_LABEL_NO_WRITE_UP (0x1)
value SYSTEM_MANDATORY_LABEL_VALID_MASK ((SYSTEM_MANDATORY_LABEL_NO_WRITE_UP | SYSTEM_MANDATORY_LABEL_NO_READ_UP | SYSTEM_MANDATORY_LABEL_NO_EXECUTE_UP))
value SYSTEM_PROCESS_TRUST_LABEL_ACE_TYPE ((0x14))
value SYSTEM_PROCESS_TRUST_LABEL_VALID_MASK (0x00ffffff)
value SYSTEM_PROCESS_TRUST_NOCONSTRAINT_MASK (0xffffffff)
value SYSTEM_RESOURCE_ATTRIBUTE_ACE_TYPE ((0x12))
value SYSTEM_SCOPED_POLICY_ID_ACE_TYPE ((0x13))
value SYSTEM_STATUS_FLAG_POWER_SAVING_ON (0x01)
value SYS_OPEN (_SYS_OPEN)
value S_ALLTHRESHOLD (2)
value S_APPLICATION_ACTIVATION_ERROR_HANDLED_BY_DIALOG (_HRESULT_TYPEDEF_(0x00270259L))
value S_ASYNCHRONOUS (MK_S_ASYNCHRONOUS)
value S_FALSE (((HRESULT)1L))
value S_IEXEC (_S_IEXEC)
value S_IFCHR (_S_IFCHR)
value S_IFDIR (_S_IFDIR)
value S_IFMT (_S_IFMT)
value S_IFREG (_S_IFREG)
value S_IREAD (_S_IREAD)
value S_IWRITE (_S_IWRITE)
value S_LEGATO (1)
value S_NORMAL (0)
value S_OK (((HRESULT)0L))
value S_PERIODVOICE (3)
value S_QUEUEEMPTY (0)
value S_SERBDNT ((-5))
value S_SERDCC ((-7))
value S_SERDDR ((-14))
value S_SERDFQ ((-13))
value S_SERDLN ((-6))
value S_SERDMD ((-10))
value S_SERDPT ((-12))
value S_SERDSH ((-11))
value S_SERDSR ((-15))
value S_SERDST ((-16))
value S_SERDTP ((-8))
value S_SERDVL ((-9))
value S_SERDVNA ((-1))
value S_SERMACT ((-3))
value S_SEROFM ((-2))
value S_SERQFUL ((-4))
value S_STACCATO (2)
value S_STORE_LAUNCHED_FOR_REMEDIATION (_HRESULT_TYPEDEF_(0x00270258L))
value S_THRESHOLD (1)
value S_WHITEVOICE (7)
value TAPE_ABSOLUTE_BLOCK (1)
value TAPE_ABSOLUTE_POSITION (0)
value TAPE_CHECK_FOR_DRIVE_PROBLEM (2)
value TAPE_DRIVE_ABSOLUTE_BLK (0x80001000)
value TAPE_DRIVE_ABS_BLK_IMMED (0x80002000)
value TAPE_DRIVE_CLEAN_REQUESTS (0x02000000)
value TAPE_DRIVE_COMPRESSION (0x00020000)
value TAPE_DRIVE_ECC (0x00010000)
value TAPE_DRIVE_EJECT_MEDIA (0x01000000)
value TAPE_DRIVE_END_OF_DATA (0x80010000)
value TAPE_DRIVE_EOT_WZ_SIZE (0x00002000)
value TAPE_DRIVE_ERASE_BOP_ONLY (0x00000040)
value TAPE_DRIVE_ERASE_IMMEDIATE (0x00000080)
value TAPE_DRIVE_ERASE_LONG (0x00000020)
value TAPE_DRIVE_ERASE_SHORT (0x00000010)
value TAPE_DRIVE_FILEMARKS (0x80040000)
value TAPE_DRIVE_FIXED (0x00000001)
value TAPE_DRIVE_FIXED_BLOCK (0x00000400)
value TAPE_DRIVE_FORMAT (0xA0000000)
value TAPE_DRIVE_FORMAT_IMMEDIATE (0xC0000000)
value TAPE_DRIVE_GET_ABSOLUTE_BLK (0x00100000)
value TAPE_DRIVE_GET_LOGICAL_BLK (0x00200000)
value TAPE_DRIVE_HIGH_FEATURES (0x80000000)
value TAPE_DRIVE_INITIATOR (0x00000004)
value TAPE_DRIVE_LOAD_UNLD_IMMED (0x80000020)
value TAPE_DRIVE_LOAD_UNLOAD (0x80000001)
value TAPE_DRIVE_LOCK_UNLK_IMMED (0x80000080)
value TAPE_DRIVE_LOCK_UNLOCK (0x80000004)
value TAPE_DRIVE_LOGICAL_BLK (0x80004000)
value TAPE_DRIVE_LOG_BLK_IMMED (0x80008000)
value TAPE_DRIVE_PADDING (0x00040000)
value TAPE_DRIVE_RELATIVE_BLKS (0x80020000)
value TAPE_DRIVE_REPORT_SMKS (0x00080000)
value TAPE_DRIVE_RESERVED_BIT (0x80000000)
value TAPE_DRIVE_REVERSE_POSITION (0x80400000)
value TAPE_DRIVE_REWIND_IMMEDIATE (0x80000008)
value TAPE_DRIVE_SELECT (0x00000002)
value TAPE_DRIVE_SEQUENTIAL_FMKS (0x80080000)
value TAPE_DRIVE_SEQUENTIAL_SMKS (0x80200000)
value TAPE_DRIVE_SETMARKS (0x80100000)
value TAPE_DRIVE_SET_BLOCK_SIZE (0x80000010)
value TAPE_DRIVE_SET_CMP_BOP_ONLY (0x04000000)
value TAPE_DRIVE_SET_COMPRESSION (0x80000200)
value TAPE_DRIVE_SET_ECC (0x80000100)
value TAPE_DRIVE_SET_EOT_WZ_SIZE (0x00400000)
value TAPE_DRIVE_SET_PADDING (0x80000400)
value TAPE_DRIVE_SET_REPORT_SMKS (0x80000800)
value TAPE_DRIVE_SPACE_IMMEDIATE (0x80800000)
value TAPE_DRIVE_TAPE_CAPACITY (0x00000100)
value TAPE_DRIVE_TAPE_REMAINING (0x00000200)
value TAPE_DRIVE_TENSION (0x80000002)
value TAPE_DRIVE_TENSION_IMMED (0x80000040)
value TAPE_DRIVE_VARIABLE_BLOCK (0x00000800)
value TAPE_DRIVE_WRITE_FILEMARKS (0x82000000)
value TAPE_DRIVE_WRITE_LONG_FMKS (0x88000000)
value TAPE_DRIVE_WRITE_MARK_IMMED (0x90000000)
value TAPE_DRIVE_WRITE_PROTECT (0x00001000)
value TAPE_DRIVE_WRITE_SETMARKS (0x81000000)
value TAPE_DRIVE_WRITE_SHORT_FMKS (0x84000000)
value TAPE_ERASE_LONG (1)
value TAPE_ERASE_SHORT (0)
value TAPE_FILEMARKS (1)
value TAPE_FIXED_PARTITIONS (0)
value TAPE_FORMAT (5)
value TAPE_INITIATOR_PARTITIONS (2)
value TAPE_LOAD (0)
value TAPE_LOCK (3)
value TAPE_LOGICAL_BLOCK (2)
value TAPE_LOGICAL_POSITION (1)
value TAPE_LONG_FILEMARKS (3)
value TAPE_PSEUDO_LOGICAL_BLOCK (3)
value TAPE_PSEUDO_LOGICAL_POSITION (2)
value TAPE_QUERY_DEVICE_ERROR_DATA (4)
value TAPE_QUERY_DRIVE_PARAMETERS (0)
value TAPE_QUERY_IO_ERROR_DATA (3)
value TAPE_QUERY_MEDIA_CAPACITY (1)
value TAPE_RESET_STATISTICS (2)
value TAPE_RETURN_ENV_INFO (1)
value TAPE_RETURN_STATISTICS (0)
value TAPE_REWIND (0)
value TAPE_SELECT_PARTITIONS (1)
value TAPE_SETMARKS (0)
value TAPE_SHORT_FILEMARKS (2)
value TAPE_SPACE_END_OF_DATA (4)
value TAPE_SPACE_FILEMARKS (6)
value TAPE_SPACE_RELATIVE_BLOCKS (5)
value TAPE_SPACE_SEQUENTIAL_FMKS (7)
value TAPE_SPACE_SEQUENTIAL_SMKS (9)
value TAPE_SPACE_SETMARKS (8)
value TAPE_TENSION (2)
value TAPE_UNLOAD (1)
value TAPE_UNLOCK (4)
value TA_BASELINE (24)
value TA_BOTTOM (8)
value TA_CENTER (6)
value TA_LEFT (0)
value TA_MASK ((TA_BASELINE+TA_CENTER+TA_UPDATECP+TA_RTLREADING))
value TA_NOUPDATECP (0)
value TA_RIGHT (2)
value TA_RTLREADING (256)
value TA_TOP (0)
value TA_UPDATECP (1)
value TBSIMP_E_BUFFER_TOO_SMALL (_HRESULT_TYPEDEF_(0x80290200L))
value TBSIMP_E_CLEANUP_FAILED (_HRESULT_TYPEDEF_(0x80290201L))
value TBSIMP_E_COMMAND_CANCELED (_HRESULT_TYPEDEF_(0x8029020BL))
value TBSIMP_E_COMMAND_FAILED (_HRESULT_TYPEDEF_(0x80290211L))
value TBSIMP_E_DUPLICATE_VHANDLE (_HRESULT_TYPEDEF_(0x80290206L))
value TBSIMP_E_HASH_BAD_KEY (_HRESULT_TYPEDEF_(0x80290205L))
value TBSIMP_E_HASH_TABLE_FULL (_HRESULT_TYPEDEF_(0x80290216L))
value TBSIMP_E_INVALID_CONTEXT_HANDLE (_HRESULT_TYPEDEF_(0x80290202L))
value TBSIMP_E_INVALID_CONTEXT_PARAM (_HRESULT_TYPEDEF_(0x80290203L))
value TBSIMP_E_INVALID_OUTPUT_POINTER (_HRESULT_TYPEDEF_(0x80290207L))
value TBSIMP_E_INVALID_PARAMETER (_HRESULT_TYPEDEF_(0x80290208L))
value TBSIMP_E_INVALID_RESOURCE (_HRESULT_TYPEDEF_(0x80290214L))
value TBSIMP_E_LIST_NOT_FOUND (_HRESULT_TYPEDEF_(0x8029020EL))
value TBSIMP_E_LIST_NO_MORE_ITEMS (_HRESULT_TYPEDEF_(0x8029020DL))
value TBSIMP_E_NOTHING_TO_UNLOAD (_HRESULT_TYPEDEF_(0x80290215L))
value TBSIMP_E_NOT_ENOUGH_SPACE (_HRESULT_TYPEDEF_(0x8029020FL))
value TBSIMP_E_NOT_ENOUGH_TPM_CONTEXTS (_HRESULT_TYPEDEF_(0x80290210L))
value TBSIMP_E_NO_EVENT_LOG (_HRESULT_TYPEDEF_(0x8029021BL))
value TBSIMP_E_OUT_OF_MEMORY (_HRESULT_TYPEDEF_(0x8029020CL))
value TBSIMP_E_PPI_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80290219L))
value TBSIMP_E_RESOURCE_EXPIRED (_HRESULT_TYPEDEF_(0x80290213L))
value TBSIMP_E_RPC_INIT_FAILED (_HRESULT_TYPEDEF_(0x80290209L))
value TBSIMP_E_SCHEDULER_NOT_RUNNING (_HRESULT_TYPEDEF_(0x8029020AL))
value TBSIMP_E_TOO_MANY_RESOURCES (_HRESULT_TYPEDEF_(0x80290218L))
value TBSIMP_E_TOO_MANY_TBS_CONTEXTS (_HRESULT_TYPEDEF_(0x80290217L))
value TBSIMP_E_TPM_ERROR (_HRESULT_TYPEDEF_(0x80290204L))
value TBSIMP_E_TPM_INCOMPATIBLE (_HRESULT_TYPEDEF_(0x8029021AL))
value TBSIMP_E_UNKNOWN_ORDINAL (_HRESULT_TYPEDEF_(0x80290212L))
value TBS_E_ACCESS_DENIED (_HRESULT_TYPEDEF_(0x80284012L))
value TBS_E_BAD_PARAMETER (_HRESULT_TYPEDEF_(0x80284002L))
value TBS_E_BUFFER_TOO_LARGE (_HRESULT_TYPEDEF_(0x8028400EL))
value TBS_E_COMMAND_CANCELED (_HRESULT_TYPEDEF_(0x8028400DL))
value TBS_E_INSUFFICIENT_BUFFER (_HRESULT_TYPEDEF_(0x80284005L))
value TBS_E_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x80284001L))
value TBS_E_INVALID_CONTEXT (_HRESULT_TYPEDEF_(0x80284004L))
value TBS_E_INVALID_CONTEXT_PARAM (_HRESULT_TYPEDEF_(0x80284007L))
value TBS_E_INVALID_OUTPUT_POINTER (_HRESULT_TYPEDEF_(0x80284003L))
value TBS_E_IOERROR (_HRESULT_TYPEDEF_(0x80284006L))
value TBS_E_NO_EVENT_LOG (_HRESULT_TYPEDEF_(0x80284011L))
value TBS_E_OWNERAUTH_NOT_FOUND (_HRESULT_TYPEDEF_(0x80284015L))
value TBS_E_PPI_FUNCTION_UNSUPPORTED (_HRESULT_TYPEDEF_(0x80284014L))
value TBS_E_PPI_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8028400CL))
value TBS_E_PROVISIONING_INCOMPLETE (_HRESULT_TYPEDEF_(0x80284016L))
value TBS_E_PROVISIONING_NOT_ALLOWED (_HRESULT_TYPEDEF_(0x80284013L))
value TBS_E_SERVICE_DISABLED (_HRESULT_TYPEDEF_(0x80284010L))
value TBS_E_SERVICE_NOT_RUNNING (_HRESULT_TYPEDEF_(0x80284008L))
value TBS_E_SERVICE_START_PENDING (_HRESULT_TYPEDEF_(0x8028400BL))
value TBS_E_TOO_MANY_RESOURCES (_HRESULT_TYPEDEF_(0x8028400AL))
value TBS_E_TOO_MANY_TBS_CONTEXTS (_HRESULT_TYPEDEF_(0x80284009L))
value TBS_E_TPM_NOT_FOUND (_HRESULT_TYPEDEF_(0x8028400FL))
value TCI_SRCCHARSET (1)
value TCI_SRCCODEPAGE (2)
value TCI_SRCFONTSIG (3)
value TCI_SRCLOCALE (0x1000)
value TCP_NODELAY (0x0001)
value TC_CP_STROKE (0x00000004)
value TC_CR_ANY (0x00000010)
value TC_DEVICEDUMP_SUBSECTION_DESC_LENGTH (16)
value TC_EA_DOUBLE (0x00000200)
value TC_GP_TRAP (2)
value TC_HARDERR (1)
value TC_IA_ABLE (0x00000400)
value TC_NONCONF_BORROW (0)
value TC_NONCONF_BORROW_PLUS (3)
value TC_NONCONF_DISCARD (2)
value TC_NONCONF_SHAPE (1)
value TC_NORMAL (0)
value TC_OP_CHARACTER (0x00000001)
value TC_OP_STROKE (0x00000002)
value TC_PUBLIC_DEVICEDUMP_CONTENT_GPLOG (0x02)
value TC_PUBLIC_DEVICEDUMP_CONTENT_GPLOG_MAX (16)
value TC_PUBLIC_DEVICEDUMP_CONTENT_SMART (0x01)
value TC_RA_ABLE (0x00002000)
value TC_RESERVED (0x00008000)
value TC_SA_CONTIN (0x00000100)
value TC_SA_DOUBLE (0x00000040)
value TC_SA_INTEGER (0x00000080)
value TC_SCROLLBLT (0x00010000)
value TC_SF_X_YINDEP (0x00000020)
value TC_SIGNAL (3)
value TC_SO_ABLE (0x00001000)
value TC_UA_ABLE (0x00000800)
value TC_VA_ABLE (0x00004000)
value TECHNOLOGY (2)
value TELEMETRY_COMMAND_SIZE (16)
value TEXTCAPS (34)
value THAI_CHARSET (222)
value THREAD_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | SYNCHRONIZE | 0xFFFF))
value THREAD_BASE_PRIORITY_IDLE ((-15))
value THREAD_BASE_PRIORITY_LOWRT (15)
value THREAD_BASE_PRIORITY_MAX (2)
value THREAD_BASE_PRIORITY_MIN ((-2))
value THREAD_DIRECT_IMPERSONATION ((0x0200))
value THREAD_DYNAMIC_CODE_ALLOW (1)
value THREAD_GET_CONTEXT ((0x0008))
value THREAD_IMPERSONATE ((0x0100))
value THREAD_MODE_BACKGROUND_BEGIN (0x00010000)
value THREAD_MODE_BACKGROUND_END (0x00020000)
value THREAD_POWER_THROTTLING_CURRENT_VERSION (1)
value THREAD_POWER_THROTTLING_EXECUTION_SPEED (0x1)
value THREAD_POWER_THROTTLING_VALID_FLAGS ((THREAD_POWER_THROTTLING_EXECUTION_SPEED))
value THREAD_PRIORITY_ABOVE_NORMAL ((THREAD_PRIORITY_HIGHEST-1))
value THREAD_PRIORITY_BELOW_NORMAL ((THREAD_PRIORITY_LOWEST+1))
value THREAD_PRIORITY_ERROR_RETURN ((MAXLONG))
value THREAD_PRIORITY_HIGHEST (THREAD_BASE_PRIORITY_MAX)
value THREAD_PRIORITY_IDLE (THREAD_BASE_PRIORITY_IDLE)
value THREAD_PRIORITY_LOWEST (THREAD_BASE_PRIORITY_MIN)
value THREAD_PRIORITY_NORMAL (0)
value THREAD_PRIORITY_TIME_CRITICAL (THREAD_BASE_PRIORITY_LOWRT)
value THREAD_PROFILING_FLAG_DISPATCH (0x00000001)
value THREAD_QUERY_INFORMATION ((0x0040))
value THREAD_QUERY_LIMITED_INFORMATION ((0x0800))
value THREAD_RESUME ((0x1000))
value THREAD_SET_CONTEXT ((0x0010))
value THREAD_SET_INFORMATION ((0x0020))
value THREAD_SET_LIMITED_INFORMATION ((0x0400))
value THREAD_SET_THREAD_TOKEN ((0x0080))
value THREAD_SUSPEND_RESUME ((0x0002))
value THREAD_TERMINATE ((0x0001))
value TH_NETDEV (0x00000001)
value TH_TAPI (0x00000002)
value TIMEFMT_ENUMPROC (TIMEFMT_ENUMPROCA)
value TIMEOUT_ASYNC (0xFFFFFFFF)
value TIMERR_BASE (96)
value TIMERR_NOCANDO ((TIMERR_BASE+1))
value TIMERR_NOERROR ((0))
value TIMERR_STRUCT ((TIMERR_BASE+33))
value TIMERV_COALESCING_MAX ((0x7FFFFFF5))
value TIMERV_COALESCING_MIN ((1))
value TIMERV_DEFAULT_COALESCING ((0))
value TIMERV_NO_COALESCING ((0xFFFFFFFF))
value TIMER_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED|SYNCHRONIZE| TIMER_QUERY_STATE|TIMER_MODIFY_STATE))
value TIMER_MODIFY_STATE (0x0002)
value TIMER_QUERY_STATE (0x0001)
value TIMESTAMP_DONT_HASH_DATA (0x00000001)
value TIMESTAMP_FAILURE_BAD_ALG (0)
value TIMESTAMP_FAILURE_BAD_FORMAT (5)
value TIMESTAMP_FAILURE_BAD_REQUEST (2)
value TIMESTAMP_FAILURE_EXTENSION_NOT_SUPPORTED (16)
value TIMESTAMP_FAILURE_INFO_NOT_AVAILABLE (17)
value TIMESTAMP_FAILURE_POLICY_NOT_SUPPORTED (15)
value TIMESTAMP_FAILURE_SYSTEM_FAILURE (25)
value TIMESTAMP_FAILURE_TIME_NOT_AVAILABLE (14)
value TIMESTAMP_INFO (((LPCSTR) 80))
value TIMESTAMP_NO_AUTH_RETRIEVAL (0x00020000)
value TIMESTAMP_REQUEST (((LPCSTR) 78))
value TIMESTAMP_RESPONSE (((LPCSTR) 79))
value TIMESTAMP_STATUS_GRANTED (0)
value TIMESTAMP_STATUS_GRANTED_WITH_MODS (1)
value TIMESTAMP_STATUS_REJECTED (2)
value TIMESTAMP_STATUS_REVOCATION_WARNING (4)
value TIMESTAMP_STATUS_REVOKED (5)
value TIMESTAMP_STATUS_WAITING (3)
value TIMESTAMP_VERIFY_CONTEXT_SIGNATURE (0x00000020)
value TIMESTAMP_VERSION (1)
value TIME_BYTES (0x0004)
value TIME_CALLBACK_EVENT_PULSE (0x0020)
value TIME_CALLBACK_EVENT_SET (0x0010)
value TIME_CALLBACK_FUNCTION (0x0000)
value TIME_KILL_SYNCHRONOUS (0x0100)
value TIME_MIDI (0x0010)
value TIME_MS (0x0001)
value TIME_NOMINUTESORSECONDS (0x00000001)
value TIME_NOSECONDS (0x00000002)
value TIME_NOTIMEMARKER (0x00000004)
value TIME_ONESHOT (0x0000)
value TIME_PERIODIC (0x0001)
value TIME_SAMPLES (0x0002)
value TIME_SMPTE (0x0008)
value TIME_TICKS (0x0020)
value TIME_UTC (1)
value TIME_VALID_OID_FLUSH_CRL (((LPCSTR)2))
value TIME_VALID_OID_FLUSH_CRL_FROM_CERT (((LPCSTR)3))
value TIME_VALID_OID_FLUSH_CTL (((LPCSTR)1))
value TIME_VALID_OID_FLUSH_FRESHEST_CRL_FROM_CERT (((LPCSTR)4))
value TIME_VALID_OID_FLUSH_FRESHEST_CRL_FROM_CRL (((LPCSTR)5))
value TIME_VALID_OID_GET_CRL (((LPCSTR)2))
value TIME_VALID_OID_GET_CRL_FROM_CERT (((LPCSTR)3))
value TIME_VALID_OID_GET_CTL (((LPCSTR)1))
value TIME_VALID_OID_GET_FRESHEST_CRL_FROM_CERT (((LPCSTR)4))
value TIME_VALID_OID_GET_FRESHEST_CRL_FROM_CRL (((LPCSTR)5))
value TIME_ZONE_ID_DAYLIGHT (2)
value TIME_ZONE_ID_INVALID (((DWORD)0xFFFFFFFF))
value TIME_ZONE_ID_STANDARD (1)
value TIME_ZONE_ID_UNKNOWN (0)
value TKF_AVAILABLE (0x00000002)
value TKF_CONFIRMHOTKEY (0x00000008)
value TKF_HOTKEYACTIVE (0x00000004)
value TKF_HOTKEYSOUND (0x00000010)
value TKF_INDICATOR (0x00000020)
value TKF_TOGGLEKEYSON (0x00000001)
value TLS_MINIMUM_AVAILABLE (64)
value TLS_OUT_OF_INDEXES (((DWORD)0xFFFFFFFF))
value TME_CANCEL (0x80000000)
value TME_HOVER (0x00000001)
value TME_LEAVE (0x00000002)
value TME_NONCLIENT (0x00000010)
value TME_QUERY (0x40000000)
value TMPF_DEVICE (0x08)
value TMPF_FIXED_PITCH (0x01)
value TMPF_TRUETYPE (0x04)
value TMPF_VECTOR (0x02)
value TMP_MAX (_CRT_INT_MAX)
value TMP_MAX_S (TMP_MAX)
value TOKEN_ACCESS_PSEUDO_HANDLE (TOKEN_ACCESS_PSEUDO_HANDLE_WIN8)
value TOKEN_ADJUST_DEFAULT ((0x0080))
value TOKEN_ADJUST_GROUPS ((0x0040))
value TOKEN_ADJUST_PRIVILEGES ((0x0020))
value TOKEN_ADJUST_SESSIONID ((0x0100))
value TOKEN_ALL_ACCESS ((TOKEN_ALL_ACCESS_P | TOKEN_ADJUST_SESSIONID ))
value TOKEN_ALL_ACCESS_P ((STANDARD_RIGHTS_REQUIRED | TOKEN_ASSIGN_PRIMARY | TOKEN_DUPLICATE | TOKEN_IMPERSONATE | TOKEN_QUERY | TOKEN_QUERY_SOURCE | TOKEN_ADJUST_PRIVILEGES | TOKEN_ADJUST_GROUPS | TOKEN_ADJUST_DEFAULT ))
value TOKEN_ASSIGN_PRIMARY ((0x0001))
value TOKEN_DUPLICATE ((0x0002))
value TOKEN_EXECUTE ((STANDARD_RIGHTS_EXECUTE))
value TOKEN_IMPERSONATE ((0x0004))
value TOKEN_MANDATORY_POLICY_NEW_PROCESS_MIN (0x2)
value TOKEN_MANDATORY_POLICY_NO_WRITE_UP (0x1)
value TOKEN_MANDATORY_POLICY_OFF (0x0)
value TOKEN_MANDATORY_POLICY_VALID_MASK ((TOKEN_MANDATORY_POLICY_NO_WRITE_UP | TOKEN_MANDATORY_POLICY_NEW_PROCESS_MIN))
value TOKEN_QUERY ((0x0008))
value TOKEN_QUERY_SOURCE ((0x0010))
value TOKEN_READ ((STANDARD_RIGHTS_READ | TOKEN_QUERY))
value TOKEN_SOURCE_LENGTH (8)
value TOKEN_TRUST_ALLOWED_MASK ((TOKEN_TRUST_CONSTRAINT_MASK | TOKEN_DUPLICATE | TOKEN_IMPERSONATE))
value TOKEN_TRUST_CONSTRAINT_MASK ((STANDARD_RIGHTS_READ | TOKEN_QUERY | TOKEN_QUERY_SOURCE ))
value TOKEN_WRITE ((STANDARD_RIGHTS_WRITE | TOKEN_ADJUST_PRIVILEGES | TOKEN_ADJUST_GROUPS | TOKEN_ADJUST_DEFAULT))
value TOUCHEVENTF_DOWN (0x0002)
value TOUCHEVENTF_INRANGE (0x0008)
value TOUCHEVENTF_MOVE (0x0001)
value TOUCHEVENTF_NOCOALESCE (0x0020)
value TOUCHEVENTF_PALM (0x0080)
value TOUCHEVENTF_PEN (0x0040)
value TOUCHEVENTF_PRIMARY (0x0010)
value TOUCHEVENTF_UP (0x0004)
value TOUCHINPUTMASKF_CONTACTAREA (0x0004)
value TOUCHINPUTMASKF_EXTRAINFO (0x0002)
value TOUCHINPUTMASKF_TIMEFROMSYSTEM (0x0001)
value TOUCHPREDICTIONPARAMETERS_DEFAULT_LATENCY (8)
value TOUCHPREDICTIONPARAMETERS_DEFAULT_SAMPLETIME (8)
value TOUCHPREDICTIONPARAMETERS_DEFAULT_USE_HW_TIMESTAMP (1)
value TOUCH_FEEDBACK_DEFAULT (0x1)
value TOUCH_FEEDBACK_INDIRECT (0x2)
value TOUCH_FEEDBACK_NONE (0x3)
value TOUCH_FLAG_NONE (0x00000000)
value TOUCH_HIT_TESTING_CLIENT (0x1)
value TOUCH_HIT_TESTING_DEFAULT (0x0)
value TOUCH_HIT_TESTING_NONE (0x2)
value TOUCH_HIT_TESTING_PROXIMITY_CLOSEST (0x0)
value TOUCH_HIT_TESTING_PROXIMITY_FARTHEST (0xFFF)
value TOUCH_MASK_CONTACTAREA (0x00000001)
value TOUCH_MASK_NONE (0x00000000)
value TOUCH_MASK_ORIENTATION (0x00000002)
value TOUCH_MASK_PRESSURE (0x00000004)
value TPC_E_INITIALIZE_FAIL (_HRESULT_TYPEDEF_(0x80040223L))
value TPC_E_INVALID_CONFIGURATION (_HRESULT_TYPEDEF_(0x80040239L))
value TPC_E_INVALID_DATA_FROM_RECOGNIZER (_HRESULT_TYPEDEF_(0x8004023AL))
value TPC_E_INVALID_INPUT_RECT (_HRESULT_TYPEDEF_(0x80040219L))
value TPC_E_INVALID_PACKET_DESCRIPTION (_HRESULT_TYPEDEF_(0x80040233L))
value TPC_E_INVALID_PROPERTY (_HRESULT_TYPEDEF_(0x80040241L))
value TPC_E_INVALID_RIGHTS (_HRESULT_TYPEDEF_(0x80040236L))
value TPC_E_INVALID_STROKE (_HRESULT_TYPEDEF_(0x80040222L))
value TPC_E_NOT_RELEVANT (_HRESULT_TYPEDEF_(0x80040232L))
value TPC_E_NO_DEFAULT_TABLET (_HRESULT_TYPEDEF_(0x80040212L))
value TPC_E_OUT_OF_ORDER_CALL (_HRESULT_TYPEDEF_(0x80040237L))
value TPC_E_QUEUE_FULL (_HRESULT_TYPEDEF_(0x80040238L))
value TPC_E_RECOGNIZER_NOT_REGISTERED (_HRESULT_TYPEDEF_(0x80040235L))
value TPC_E_UNKNOWN_PROPERTY (_HRESULT_TYPEDEF_(0x8004021BL))
value TPC_S_INTERRUPTED (_HRESULT_TYPEDEF_(0x00040253L))
value TPC_S_NO_DATA_TO_PROCESS (_HRESULT_TYPEDEF_(0x00040254L))
value TPC_S_TRUNCATED (_HRESULT_TYPEDEF_(0x00040252L))
value TPMAPI_E_ACCESS_DENIED (_HRESULT_TYPEDEF_(0x80290108L))
value TPMAPI_E_AUTHORIZATION_FAILED (_HRESULT_TYPEDEF_(0x80290109L))
value TPMAPI_E_AUTHORIZATION_REVOKED (_HRESULT_TYPEDEF_(0x80290126L))
value TPMAPI_E_AUTHORIZING_KEY_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80290128L))
value TPMAPI_E_BUFFER_TOO_SMALL (_HRESULT_TYPEDEF_(0x80290106L))
value TPMAPI_E_EMPTY_TCG_LOG (_HRESULT_TYPEDEF_(0x8029011AL))
value TPMAPI_E_ENCRYPTION_FAILED (_HRESULT_TYPEDEF_(0x80290110L))
value TPMAPI_E_ENDORSEMENT_AUTH_NOT_NULL (_HRESULT_TYPEDEF_(0x80290125L))
value TPMAPI_E_FIPS_RNG_CHECK_FAILED (_HRESULT_TYPEDEF_(0x80290119L))
value TPMAPI_E_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x80290107L))
value TPMAPI_E_INVALID_AUTHORIZATION_SIGNATURE (_HRESULT_TYPEDEF_(0x80290129L))
value TPMAPI_E_INVALID_CONTEXT_HANDLE (_HRESULT_TYPEDEF_(0x8029010AL))
value TPMAPI_E_INVALID_CONTEXT_PARAMS (_HRESULT_TYPEDEF_(0x80290115L))
value TPMAPI_E_INVALID_DELEGATE_BLOB (_HRESULT_TYPEDEF_(0x80290114L))
value TPMAPI_E_INVALID_ENCODING (_HRESULT_TYPEDEF_(0x8029010EL))
value TPMAPI_E_INVALID_KEY_BLOB (_HRESULT_TYPEDEF_(0x80290116L))
value TPMAPI_E_INVALID_KEY_PARAMS (_HRESULT_TYPEDEF_(0x80290111L))
value TPMAPI_E_INVALID_KEY_SIZE (_HRESULT_TYPEDEF_(0x8029010FL))
value TPMAPI_E_INVALID_MIGRATION_AUTHORIZATION_BLOB (_HRESULT_TYPEDEF_(0x80290112L))
value TPMAPI_E_INVALID_OUTPUT_POINTER (_HRESULT_TYPEDEF_(0x80290103L))
value TPMAPI_E_INVALID_OWNER_AUTH (_HRESULT_TYPEDEF_(0x80290118L))
value TPMAPI_E_INVALID_PARAMETER (_HRESULT_TYPEDEF_(0x80290104L))
value TPMAPI_E_INVALID_PCR_DATA (_HRESULT_TYPEDEF_(0x80290117L))
value TPMAPI_E_INVALID_PCR_INDEX (_HRESULT_TYPEDEF_(0x80290113L))
value TPMAPI_E_INVALID_POLICYAUTH_BLOB_TYPE (_HRESULT_TYPEDEF_(0x8029012EL))
value TPMAPI_E_INVALID_STATE (_HRESULT_TYPEDEF_(0x80290100L))
value TPMAPI_E_INVALID_TCG_LOG_ENTRY (_HRESULT_TYPEDEF_(0x8029011BL))
value TPMAPI_E_INVALID_TPM_VERSION (_HRESULT_TYPEDEF_(0x8029012DL))
value TPMAPI_E_MALFORMED_AUTHORIZATION_KEY (_HRESULT_TYPEDEF_(0x80290127L))
value TPMAPI_E_MALFORMED_AUTHORIZATION_OTHER (_HRESULT_TYPEDEF_(0x8029012BL))
value TPMAPI_E_MALFORMED_AUTHORIZATION_POLICY (_HRESULT_TYPEDEF_(0x8029012AL))
value TPMAPI_E_MESSAGE_TOO_LARGE (_HRESULT_TYPEDEF_(0x8029010DL))
value TPMAPI_E_NOT_ENOUGH_DATA (_HRESULT_TYPEDEF_(0x80290101L))
value TPMAPI_E_NO_AUTHORIZATION_CHAIN_FOUND (_HRESULT_TYPEDEF_(0x80290122L))
value TPMAPI_E_NV_BITS_NOT_DEFINED (_HRESULT_TYPEDEF_(0x8029011FL))
value TPMAPI_E_NV_BITS_NOT_READY (_HRESULT_TYPEDEF_(0x80290120L))
value TPMAPI_E_OUT_OF_MEMORY (_HRESULT_TYPEDEF_(0x80290105L))
value TPMAPI_E_OWNER_AUTH_NOT_NULL (_HRESULT_TYPEDEF_(0x80290124L))
value TPMAPI_E_POLICY_DENIES_OPERATION (_HRESULT_TYPEDEF_(0x8029011EL))
value TPMAPI_E_SEALING_KEY_CHANGED (_HRESULT_TYPEDEF_(0x8029012CL))
value TPMAPI_E_SEALING_KEY_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x80290121L))
value TPMAPI_E_SVN_COUNTER_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x80290123L))
value TPMAPI_E_TBS_COMMUNICATION_ERROR (_HRESULT_TYPEDEF_(0x8029010BL))
value TPMAPI_E_TCG_INVALID_DIGEST_ENTRY (_HRESULT_TYPEDEF_(0x8029011DL))
value TPMAPI_E_TCG_SEPARATOR_ABSENT (_HRESULT_TYPEDEF_(0x8029011CL))
value TPMAPI_E_TOO_MUCH_DATA (_HRESULT_TYPEDEF_(0x80290102L))
value TPMAPI_E_TPM_COMMAND_ERROR (_HRESULT_TYPEDEF_(0x8029010CL))
value TPM_BOTTOMALIGN (0x0020L)
value TPM_CENTERALIGN (0x0004L)
value TPM_E_AREA_LOCKED (_HRESULT_TYPEDEF_(0x8028003CL))
value TPM_E_ATTESTATION_CHALLENGE_NOT_SET (_HRESULT_TYPEDEF_(0x80290412L))
value TPM_E_AUDITFAILURE (_HRESULT_TYPEDEF_(0x80280004L))
value TPM_E_AUDITFAIL_SUCCESSFUL (_HRESULT_TYPEDEF_(0x80280031L))
value TPM_E_AUDITFAIL_UNSUCCESSFUL (_HRESULT_TYPEDEF_(0x80280030L))
value TPM_E_AUTHFAIL (_HRESULT_TYPEDEF_(0x80280001L))
value TPM_E_AUTH_CONFLICT (_HRESULT_TYPEDEF_(0x8028003BL))
value TPM_E_BADCONTEXT (_HRESULT_TYPEDEF_(0x8028005AL))
value TPM_E_BADINDEX (_HRESULT_TYPEDEF_(0x80280002L))
value TPM_E_BADTAG (_HRESULT_TYPEDEF_(0x8028001EL))
value TPM_E_BAD_ATTRIBUTES (_HRESULT_TYPEDEF_(0x80280042L))
value TPM_E_BAD_COUNTER (_HRESULT_TYPEDEF_(0x80280045L))
value TPM_E_BAD_DATASIZE (_HRESULT_TYPEDEF_(0x8028002BL))
value TPM_E_BAD_DELEGATE (_HRESULT_TYPEDEF_(0x80280059L))
value TPM_E_BAD_HANDLE (_HRESULT_TYPEDEF_(0x80280058L))
value TPM_E_BAD_KEY_PROPERTY (_HRESULT_TYPEDEF_(0x80280028L))
value TPM_E_BAD_LOCALITY (_HRESULT_TYPEDEF_(0x8028003DL))
value TPM_E_BAD_MIGRATION (_HRESULT_TYPEDEF_(0x80280029L))
value TPM_E_BAD_MODE (_HRESULT_TYPEDEF_(0x8028002CL))
value TPM_E_BAD_ORDINAL (_HRESULT_TYPEDEF_(0x8028000AL))
value TPM_E_BAD_PARAMETER (_HRESULT_TYPEDEF_(0x80280003L))
value TPM_E_BAD_PARAM_SIZE (_HRESULT_TYPEDEF_(0x80280019L))
value TPM_E_BAD_PRESENCE (_HRESULT_TYPEDEF_(0x8028002DL))
value TPM_E_BAD_SCHEME (_HRESULT_TYPEDEF_(0x8028002AL))
value TPM_E_BAD_SIGNATURE (_HRESULT_TYPEDEF_(0x80280062L))
value TPM_E_BAD_TYPE (_HRESULT_TYPEDEF_(0x80280034L))
value TPM_E_BAD_VERSION (_HRESULT_TYPEDEF_(0x8028002EL))
value TPM_E_BUFFER_LENGTH_MISMATCH (_HRESULT_TYPEDEF_(0x8029041EL))
value TPM_E_CLAIM_TYPE_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8029041CL))
value TPM_E_CLEAR_DISABLED (_HRESULT_TYPEDEF_(0x80280005L))
value TPM_E_COMMAND_BLOCKED (_HRESULT_TYPEDEF_(0x80280400L))
value TPM_E_CONTEXT_GAP (_HRESULT_TYPEDEF_(0x80280047L))
value TPM_E_DAA_ISSUER_SETTINGS (_HRESULT_TYPEDEF_(0x80280053L))
value TPM_E_DAA_ISSUER_VALIDITY (_HRESULT_TYPEDEF_(0x80280056L))
value TPM_E_DAA_RESOURCES (_HRESULT_TYPEDEF_(0x80280050L))
value TPM_E_DAA_STAGE (_HRESULT_TYPEDEF_(0x80280055L))
value TPM_E_DAA_TPM_SETTINGS (_HRESULT_TYPEDEF_(0x80280054L))
value TPM_E_DAA_WRONG_W (_HRESULT_TYPEDEF_(0x80280057L))
value TPM_E_DEACTIVATED (_HRESULT_TYPEDEF_(0x80280006L))
value TPM_E_DECRYPT_ERROR (_HRESULT_TYPEDEF_(0x80280021L))
value TPM_E_DEFEND_LOCK_RUNNING (_HRESULT_TYPEDEF_(0x80280803L))
value TPM_E_DELEGATE_ADMIN (_HRESULT_TYPEDEF_(0x8028004DL))
value TPM_E_DELEGATE_FAMILY (_HRESULT_TYPEDEF_(0x8028004CL))
value TPM_E_DELEGATE_LOCK (_HRESULT_TYPEDEF_(0x8028004BL))
value TPM_E_DISABLED (_HRESULT_TYPEDEF_(0x80280007L))
value TPM_E_DISABLED_CMD (_HRESULT_TYPEDEF_(0x80280008L))
value TPM_E_DOING_SELFTEST (_HRESULT_TYPEDEF_(0x80280802L))
value TPM_E_DUPLICATE_VHANDLE (_HRESULT_TYPEDEF_(0x80280402L))
value TPM_E_EMBEDDED_COMMAND_BLOCKED (_HRESULT_TYPEDEF_(0x80280403L))
value TPM_E_EMBEDDED_COMMAND_UNSUPPORTED (_HRESULT_TYPEDEF_(0x80280404L))
value TPM_E_ENCRYPT_ERROR (_HRESULT_TYPEDEF_(0x80280020L))
value TPM_E_ERROR_MASK (_HRESULT_TYPEDEF_(0x80280000L))
value TPM_E_FAIL (_HRESULT_TYPEDEF_(0x80280009L))
value TPM_E_FAILEDSELFTEST (_HRESULT_TYPEDEF_(0x8028001CL))
value TPM_E_FAMILYCOUNT (_HRESULT_TYPEDEF_(0x80280040L))
value TPM_E_INAPPROPRIATE_ENC (_HRESULT_TYPEDEF_(0x8028000EL))
value TPM_E_INAPPROPRIATE_SIG (_HRESULT_TYPEDEF_(0x80280027L))
value TPM_E_INSTALL_DISABLED (_HRESULT_TYPEDEF_(0x8028000BL))
value TPM_E_INVALID_AUTHHANDLE (_HRESULT_TYPEDEF_(0x80280022L))
value TPM_E_INVALID_FAMILY (_HRESULT_TYPEDEF_(0x80280037L))
value TPM_E_INVALID_HANDLE (_HRESULT_TYPEDEF_(0x80280401L))
value TPM_E_INVALID_KEYHANDLE (_HRESULT_TYPEDEF_(0x8028000CL))
value TPM_E_INVALID_KEYUSAGE (_HRESULT_TYPEDEF_(0x80280024L))
value TPM_E_INVALID_OWNER_AUTH (_HRESULT_TYPEDEF_(0x80290601L))
value TPM_E_INVALID_PCR_INFO (_HRESULT_TYPEDEF_(0x80280010L))
value TPM_E_INVALID_POSTINIT (_HRESULT_TYPEDEF_(0x80280026L))
value TPM_E_INVALID_RESOURCE (_HRESULT_TYPEDEF_(0x80280035L))
value TPM_E_INVALID_STRUCTURE (_HRESULT_TYPEDEF_(0x80280043L))
value TPM_E_IOERROR (_HRESULT_TYPEDEF_(0x8028001FL))
value TPM_E_KEYNOTFOUND (_HRESULT_TYPEDEF_(0x8028000DL))
value TPM_E_KEY_ALREADY_FINALIZED (_HRESULT_TYPEDEF_(0x80290414L))
value TPM_E_KEY_NOTSUPPORTED (_HRESULT_TYPEDEF_(0x8028003AL))
value TPM_E_KEY_NOT_AUTHENTICATED (_HRESULT_TYPEDEF_(0x80290418L))
value TPM_E_KEY_NOT_FINALIZED (_HRESULT_TYPEDEF_(0x80290411L))
value TPM_E_KEY_NOT_LOADED (_HRESULT_TYPEDEF_(0x8029040FL))
value TPM_E_KEY_NOT_SIGNING_KEY (_HRESULT_TYPEDEF_(0x8029041AL))
value TPM_E_KEY_OWNER_CONTROL (_HRESULT_TYPEDEF_(0x80280044L))
value TPM_E_KEY_USAGE_POLICY_INVALID (_HRESULT_TYPEDEF_(0x80290416L))
value TPM_E_KEY_USAGE_POLICY_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80290415L))
value TPM_E_LOCKED_OUT (_HRESULT_TYPEDEF_(0x8029041BL))
value TPM_E_MAXNVWRITES (_HRESULT_TYPEDEF_(0x80280048L))
value TPM_E_MA_AUTHORITY (_HRESULT_TYPEDEF_(0x8028005FL))
value TPM_E_MA_DESTINATION (_HRESULT_TYPEDEF_(0x8028005DL))
value TPM_E_MA_SOURCE (_HRESULT_TYPEDEF_(0x8028005EL))
value TPM_E_MA_TICKET_SIGNATURE (_HRESULT_TYPEDEF_(0x8028005CL))
value TPM_E_MIGRATEFAIL (_HRESULT_TYPEDEF_(0x8028000FL))
value TPM_E_NEEDS_SELFTEST (_HRESULT_TYPEDEF_(0x80280801L))
value TPM_E_NOCONTEXTSPACE (_HRESULT_TYPEDEF_(0x80280063L))
value TPM_E_NOOPERATOR (_HRESULT_TYPEDEF_(0x80280049L))
value TPM_E_NOSPACE (_HRESULT_TYPEDEF_(0x80280011L))
value TPM_E_NOSRK (_HRESULT_TYPEDEF_(0x80280012L))
value TPM_E_NOTFIPS (_HRESULT_TYPEDEF_(0x80280036L))
value TPM_E_NOTLOCAL (_HRESULT_TYPEDEF_(0x80280033L))
value TPM_E_NOTRESETABLE (_HRESULT_TYPEDEF_(0x80280032L))
value TPM_E_NOTSEALED_BLOB (_HRESULT_TYPEDEF_(0x80280013L))
value TPM_E_NOT_FULLWRITE (_HRESULT_TYPEDEF_(0x80280046L))
value TPM_E_NOT_PCR_BOUND (_HRESULT_TYPEDEF_(0x80290413L))
value TPM_E_NO_ENDORSEMENT (_HRESULT_TYPEDEF_(0x80280023L))
value TPM_E_NO_KEY_CERTIFICATION (_HRESULT_TYPEDEF_(0x80290410L))
value TPM_E_NO_NV_PERMISSION (_HRESULT_TYPEDEF_(0x80280038L))
value TPM_E_NO_WRAP_TRANSPORT (_HRESULT_TYPEDEF_(0x8028002FL))
value TPM_E_OWNER_CONTROL (_HRESULT_TYPEDEF_(0x8028004FL))
value TPM_E_OWNER_SET (_HRESULT_TYPEDEF_(0x80280014L))
value TPM_E_PCP_AUTHENTICATION_FAILED (_HRESULT_TYPEDEF_(0x80290408L))
value TPM_E_PCP_AUTHENTICATION_IGNORED (_HRESULT_TYPEDEF_(0x80290409L))
value TPM_E_PCP_BUFFER_TOO_SMALL (_HRESULT_TYPEDEF_(0x80290406L))
value TPM_E_PCP_DEVICE_NOT_READY (_HRESULT_TYPEDEF_(0x80290401L))
value TPM_E_PCP_ERROR_MASK (_HRESULT_TYPEDEF_(0x80290400L))
value TPM_E_PCP_FLAG_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80290404L))
value TPM_E_PCP_IFX_RSA_KEY_CREATION_BLOCKED (_HRESULT_TYPEDEF_(0x8029041FL))
value TPM_E_PCP_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x80290407L))
value TPM_E_PCP_INVALID_HANDLE (_HRESULT_TYPEDEF_(0x80290402L))
value TPM_E_PCP_INVALID_PARAMETER (_HRESULT_TYPEDEF_(0x80290403L))
value TPM_E_PCP_KEY_HANDLE_INVALIDATED (_HRESULT_TYPEDEF_(0x80290422L))
value TPM_E_PCP_KEY_NOT_AIK (_HRESULT_TYPEDEF_(0x80290419L))
value TPM_E_PCP_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80290405L))
value TPM_E_PCP_PLATFORM_CLAIM_MAY_BE_OUTDATED (_HRESULT_TYPEDEF_(0x40290424L))
value TPM_E_PCP_PLATFORM_CLAIM_OUTDATED (_HRESULT_TYPEDEF_(0x40290425L))
value TPM_E_PCP_PLATFORM_CLAIM_REBOOT (_HRESULT_TYPEDEF_(0x40290426L))
value TPM_E_PCP_POLICY_NOT_FOUND (_HRESULT_TYPEDEF_(0x8029040AL))
value TPM_E_PCP_PROFILE_NOT_FOUND (_HRESULT_TYPEDEF_(0x8029040BL))
value TPM_E_PCP_RAW_POLICY_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80290421L))
value TPM_E_PCP_TICKET_MISSING (_HRESULT_TYPEDEF_(0x80290420L))
value TPM_E_PCP_UNSUPPORTED_PSS_SALT (_HRESULT_TYPEDEF_(0x40290423L))
value TPM_E_PCP_VALIDATION_FAILED (_HRESULT_TYPEDEF_(0x8029040CL))
value TPM_E_PCP_WRONG_PARENT (_HRESULT_TYPEDEF_(0x8029040EL))
value TPM_E_PERMANENTEK (_HRESULT_TYPEDEF_(0x80280061L))
value TPM_E_PER_NOWRITE (_HRESULT_TYPEDEF_(0x8028003FL))
value TPM_E_PPI_ACPI_FAILURE (_HRESULT_TYPEDEF_(0x80290300L))
value TPM_E_PPI_BIOS_FAILURE (_HRESULT_TYPEDEF_(0x80290302L))
value TPM_E_PPI_BLOCKED_IN_BIOS (_HRESULT_TYPEDEF_(0x80290304L))
value TPM_E_PPI_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x80290303L))
value TPM_E_PPI_USER_ABORT (_HRESULT_TYPEDEF_(0x80290301L))
value TPM_E_PROVISIONING_INCOMPLETE (_HRESULT_TYPEDEF_(0x80290600L))
value TPM_E_READ_ONLY (_HRESULT_TYPEDEF_(0x8028003EL))
value TPM_E_REQUIRES_SIGN (_HRESULT_TYPEDEF_(0x80280039L))
value TPM_E_RESOURCEMISSING (_HRESULT_TYPEDEF_(0x8028004AL))
value TPM_E_RESOURCES (_HRESULT_TYPEDEF_(0x80280015L))
value TPM_E_RETRY (_HRESULT_TYPEDEF_(0x80280800L))
value TPM_E_SHA_ERROR (_HRESULT_TYPEDEF_(0x8028001BL))
value TPM_E_SHA_THREAD (_HRESULT_TYPEDEF_(0x8028001AL))
value TPM_E_SHORTRANDOM (_HRESULT_TYPEDEF_(0x80280016L))
value TPM_E_SIZE (_HRESULT_TYPEDEF_(0x80280017L))
value TPM_E_SOFT_KEY_ERROR (_HRESULT_TYPEDEF_(0x80290417L))
value TPM_E_TOOMANYCONTEXTS (_HRESULT_TYPEDEF_(0x8028005BL))
value TPM_E_TOO_MUCH_DATA (_HRESULT_TYPEDEF_(0x80290602L))
value TPM_E_TPM_GENERATED_EPS (_HRESULT_TYPEDEF_(0x80290603L))
value TPM_E_TRANSPORT_NOTEXCLUSIVE (_HRESULT_TYPEDEF_(0x8028004EL))
value TPM_E_VERSION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x8029041DL))
value TPM_E_WRITE_LOCKED (_HRESULT_TYPEDEF_(0x80280041L))
value TPM_E_WRONGPCRVAL (_HRESULT_TYPEDEF_(0x80280018L))
value TPM_E_WRONG_ENTITYTYPE (_HRESULT_TYPEDEF_(0x80280025L))
value TPM_E_ZERO_EXHAUST_ENABLED (_HRESULT_TYPEDEF_(0x80290500L))
value TPM_HORIZONTAL (0x0000L)
value TPM_HORNEGANIMATION (0x0800L)
value TPM_HORPOSANIMATION (0x0400L)
value TPM_LAYOUTRTL (0x8000L)
value TPM_LEFTALIGN (0x0000L)
value TPM_LEFTBUTTON (0x0000L)
value TPM_NOANIMATION (0x4000L)
value TPM_NONOTIFY (0x0080L)
value TPM_RECURSE (0x0001L)
value TPM_RETURNCMD (0x0100L)
value TPM_RIGHTALIGN (0x0008L)
value TPM_RIGHTBUTTON (0x0002L)
value TPM_TOPALIGN (0x0000L)
value TPM_VCENTERALIGN (0x0010L)
value TPM_VERNEGANIMATION (0x2000L)
value TPM_VERPOSANIMATION (0x1000L)
value TPM_VERTICAL (0x0040L)
value TPM_WORKAREA (0x10000L)
value TRANSACTIONMANAGER_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | TRANSACTIONMANAGER_GENERIC_READ | TRANSACTIONMANAGER_GENERIC_WRITE | TRANSACTIONMANAGER_GENERIC_EXECUTE | TRANSACTIONMANAGER_BIND_TRANSACTION))
value TRANSACTIONMANAGER_BIND_TRANSACTION (( 0x0020 ))
value TRANSACTIONMANAGER_CREATE_RM (( 0x0010 ))
value TRANSACTIONMANAGER_GENERIC_EXECUTE ((STANDARD_RIGHTS_EXECUTE))
value TRANSACTIONMANAGER_GENERIC_READ ((STANDARD_RIGHTS_READ | TRANSACTIONMANAGER_QUERY_INFORMATION))
value TRANSACTIONMANAGER_GENERIC_WRITE ((STANDARD_RIGHTS_WRITE | TRANSACTIONMANAGER_SET_INFORMATION | TRANSACTIONMANAGER_RECOVER | TRANSACTIONMANAGER_RENAME | TRANSACTIONMANAGER_CREATE_RM))
value TRANSACTIONMANAGER_QUERY_INFORMATION (( 0x0001 ))
value TRANSACTIONMANAGER_RECOVER (( 0x0004 ))
value TRANSACTIONMANAGER_RENAME (( 0x0008 ))
value TRANSACTIONMANAGER_SET_INFORMATION (( 0x0002 ))
value TRANSACTION_ALL_ACCESS ((STANDARD_RIGHTS_REQUIRED | TRANSACTION_GENERIC_READ | TRANSACTION_GENERIC_WRITE | TRANSACTION_GENERIC_EXECUTE))
value TRANSACTION_COMMIT (( 0x0008 ))
value TRANSACTION_DO_NOT_PROMOTE (0x00000001)
value TRANSACTION_ENLIST (( 0x0004 ))
value TRANSACTION_GENERIC_EXECUTE ((STANDARD_RIGHTS_EXECUTE | TRANSACTION_COMMIT | TRANSACTION_ROLLBACK | SYNCHRONIZE))
value TRANSACTION_GENERIC_READ ((STANDARD_RIGHTS_READ | TRANSACTION_QUERY_INFORMATION | SYNCHRONIZE))
value TRANSACTION_GENERIC_WRITE ((STANDARD_RIGHTS_WRITE | TRANSACTION_SET_INFORMATION | TRANSACTION_COMMIT | TRANSACTION_ENLIST | TRANSACTION_ROLLBACK | TRANSACTION_PROPAGATE | SYNCHRONIZE))
value TRANSACTION_MANAGER_COMMIT_DEFAULT (0x00000000)
value TRANSACTION_MANAGER_COMMIT_LOWEST (0x00000008)
value TRANSACTION_MANAGER_COMMIT_SYSTEM_HIVES (0x00000004)
value TRANSACTION_MANAGER_COMMIT_SYSTEM_VOLUME (0x00000002)
value TRANSACTION_MANAGER_CORRUPT_FOR_PROGRESS (0x00000020)
value TRANSACTION_MANAGER_CORRUPT_FOR_RECOVERY (0x00000010)
value TRANSACTION_MANAGER_MAXIMUM_OPTION (0x0000003F)
value TRANSACTION_MANAGER_VOLATILE (0x00000001)
value TRANSACTION_MAXIMUM_OPTION (0x00000001)
value TRANSACTION_NOTIFICATION_TM_ONLINE_FLAG_IS_CLUSTERED (0x1)
value TRANSACTION_NOTIFY_COMMIT (0x00000004)
value TRANSACTION_NOTIFY_COMMIT_COMPLETE (0x00000040)
value TRANSACTION_NOTIFY_COMMIT_FINALIZE (0x40000000)
value TRANSACTION_NOTIFY_COMMIT_REQUEST (0x04000000)
value TRANSACTION_NOTIFY_DELEGATE_COMMIT (0x00000400)
value TRANSACTION_NOTIFY_ENLIST_MASK (0x00040000)
value TRANSACTION_NOTIFY_ENLIST_PREPREPARE (0x00001000)
value TRANSACTION_NOTIFY_INDOUBT (0x00004000)
value TRANSACTION_NOTIFY_LAST_RECOVER (0x00002000)
value TRANSACTION_NOTIFY_MARSHAL (0x00020000)
value TRANSACTION_NOTIFY_MASK (0x3FFFFFFF)
value TRANSACTION_NOTIFY_PREPARE (0x00000002)
value TRANSACTION_NOTIFY_PREPARE_COMPLETE (0x00000020)
value TRANSACTION_NOTIFY_PREPREPARE (0x00000001)
value TRANSACTION_NOTIFY_PREPREPARE_COMPLETE (0x00000010)
value TRANSACTION_NOTIFY_PROMOTE (0x08000000)
value TRANSACTION_NOTIFY_PROMOTE_NEW (0x10000000)
value TRANSACTION_NOTIFY_PROPAGATE_PULL (0x00008000)
value TRANSACTION_NOTIFY_PROPAGATE_PUSH (0x00010000)
value TRANSACTION_NOTIFY_RECOVER (0x00000100)
value TRANSACTION_NOTIFY_RECOVER_QUERY (0x00000800)
value TRANSACTION_NOTIFY_REQUEST_OUTCOME (0x20000000)
value TRANSACTION_NOTIFY_RM_DISCONNECTED (0x01000000)
value TRANSACTION_NOTIFY_ROLLBACK (0x00000008)
value TRANSACTION_NOTIFY_ROLLBACK_COMPLETE (0x00000080)
value TRANSACTION_NOTIFY_SINGLE_PHASE_COMMIT (0x00000200)
value TRANSACTION_NOTIFY_TM_ONLINE (0x02000000)
value TRANSACTION_PROPAGATE (( 0x0020 ))
value TRANSACTION_QUERY_INFORMATION (( 0x0001 ))
value TRANSACTION_RESOURCE_MANAGER_RIGHTS ((TRANSACTION_GENERIC_READ | STANDARD_RIGHTS_WRITE | TRANSACTION_SET_INFORMATION | TRANSACTION_ENLIST | TRANSACTION_ROLLBACK | TRANSACTION_PROPAGATE | SYNCHRONIZE))
value TRANSACTION_ROLLBACK (( 0x0010 ))
value TRANSACTION_SET_INFORMATION (( 0x0002 ))
value TRANSFORM_CTM (4107)
value TRANSPARENT (1)
value TRANSPORT_TYPE_CN (0x01)
value TRANSPORT_TYPE_DG (0x02)
value TRANSPORT_TYPE_LPC (0x04)
value TRANSPORT_TYPE_WMSG (0x08)
value TREE_CONNECT_ATTRIBUTE_GLOBAL (0x00000004)
value TREE_CONNECT_ATTRIBUTE_INTEGRITY (0x00008000)
value TREE_CONNECT_ATTRIBUTE_PINNED (0x00000002)
value TREE_CONNECT_ATTRIBUTE_PRIVACY (0x00004000)
value TRUE (1)
value TRUETYPE_FONTTYPE (0x0004)
value TRUNCATE_EXISTING (5)
value TRUST_E_ACTION_UNKNOWN (_HRESULT_TYPEDEF_(0x800B0002L))
value TRUST_E_BAD_DIGEST (_HRESULT_TYPEDEF_(0x80096010L))
value TRUST_E_BASIC_CONSTRAINTS (_HRESULT_TYPEDEF_(0x80096019L))
value TRUST_E_CERT_SIGNATURE (_HRESULT_TYPEDEF_(0x80096004L))
value TRUST_E_COUNTER_SIGNER (_HRESULT_TYPEDEF_(0x80096003L))
value TRUST_E_EXPLICIT_DISTRUST (_HRESULT_TYPEDEF_(0x800B0111L))
value TRUST_E_FAIL (_HRESULT_TYPEDEF_(0x800B010BL))
value TRUST_E_FINANCIAL_CRITERIA (_HRESULT_TYPEDEF_(0x8009601EL))
value TRUST_E_MALFORMED_SIGNATURE (_HRESULT_TYPEDEF_(0x80096011L))
value TRUST_E_NOSIGNATURE (_HRESULT_TYPEDEF_(0x800B0100L))
value TRUST_E_NO_SIGNER_CERT (_HRESULT_TYPEDEF_(0x80096002L))
value TRUST_E_PROVIDER_UNKNOWN (_HRESULT_TYPEDEF_(0x800B0001L))
value TRUST_E_SUBJECT_FORM_UNKNOWN (_HRESULT_TYPEDEF_(0x800B0003L))
value TRUST_E_SUBJECT_NOT_TRUSTED (_HRESULT_TYPEDEF_(0x800B0004L))
value TRUST_E_SYSTEM_ERROR (_HRESULT_TYPEDEF_(0x80096001L))
value TRUST_E_TIME_STAMP (_HRESULT_TYPEDEF_(0x80096005L))
value TRUST_PROTECTED_FILTER_ACE_FLAG ((0x40))
value TRY_AGAIN (WSATRY_AGAIN)
value TT_AVAILABLE (0x0001)
value TT_ENABLED (0x0002)
value TT_OPENTYPE_FONTTYPE (0x20000)
value TT_POLYGON_TYPE (24)
value TT_PRIM_CSPLINE (3)
value TT_PRIM_LINE (1)
value TT_PRIM_QSPLINE (2)
value TURKISH_CHARSET (162)
value TWF_FINETOUCH ((0x00000001))
value TWF_WANTPALM ((0x00000002))
value TWOSTOPBITS (2)
value TXFS_LIST_TRANSACTION_LOCKED_FILES_ENTRY_FLAG_CREATED (0x00000001)
value TXFS_LIST_TRANSACTION_LOCKED_FILES_ENTRY_FLAG_DELETED (0x00000002)
value TXFS_LOGGING_MODE_FULL ((0x0002))
value TXFS_LOGGING_MODE_SIMPLE ((0x0001))
value TXFS_MODIFY_RM_VALID_FLAGS ((TXFS_RM_FLAG_LOGGING_MODE | TXFS_RM_FLAG_RENAME_RM | TXFS_RM_FLAG_LOG_CONTAINER_COUNT_MAX | TXFS_RM_FLAG_LOG_CONTAINER_COUNT_MIN | TXFS_RM_FLAG_LOG_GROWTH_INCREMENT_NUM_CONTAINERS | TXFS_RM_FLAG_LOG_GROWTH_INCREMENT_PERCENT | TXFS_RM_FLAG_LOG_AUTO_SHRINK_PERCENTAGE | TXFS_RM_FLAG_LOG_NO_CONTAINER_COUNT_MAX | TXFS_RM_FLAG_LOG_NO_CONTAINER_COUNT_MIN | TXFS_RM_FLAG_SHRINK_LOG | TXFS_RM_FLAG_GROW_LOG | TXFS_RM_FLAG_ENFORCE_MINIMUM_SIZE | TXFS_RM_FLAG_PRESERVE_CHANGES | TXFS_RM_FLAG_RESET_RM_AT_NEXT_START | TXFS_RM_FLAG_DO_NOT_RESET_RM_AT_NEXT_START | TXFS_RM_FLAG_PREFER_CONSISTENCY | TXFS_RM_FLAG_PREFER_AVAILABILITY))
value TXFS_QUERY_RM_INFORMATION_VALID_FLAGS ((TXFS_RM_FLAG_LOG_GROWTH_INCREMENT_NUM_CONTAINERS | TXFS_RM_FLAG_LOG_GROWTH_INCREMENT_PERCENT | TXFS_RM_FLAG_LOG_NO_CONTAINER_COUNT_MAX | TXFS_RM_FLAG_LOG_NO_CONTAINER_COUNT_MIN | TXFS_RM_FLAG_RESET_RM_AT_NEXT_START | TXFS_RM_FLAG_DO_NOT_RESET_RM_AT_NEXT_START | TXFS_RM_FLAG_PREFER_CONSISTENCY | TXFS_RM_FLAG_PREFER_AVAILABILITY))
value TXFS_RM_FLAG_DO_NOT_RESET_RM_AT_NEXT_START (0x00008000)
value TXFS_RM_FLAG_ENFORCE_MINIMUM_SIZE (0x00001000)
value TXFS_RM_FLAG_GROW_LOG (0x00000400)
value TXFS_RM_FLAG_LOGGING_MODE (0x00000001)
value TXFS_RM_FLAG_LOG_AUTO_SHRINK_PERCENTAGE (0x00000040)
value TXFS_RM_FLAG_LOG_CONTAINER_COUNT_MAX (0x00000004)
value TXFS_RM_FLAG_LOG_CONTAINER_COUNT_MIN (0x00000008)
value TXFS_RM_FLAG_LOG_GROWTH_INCREMENT_NUM_CONTAINERS (0x00000010)
value TXFS_RM_FLAG_LOG_GROWTH_INCREMENT_PERCENT (0x00000020)
value TXFS_RM_FLAG_LOG_NO_CONTAINER_COUNT_MAX (0x00000080)
value TXFS_RM_FLAG_LOG_NO_CONTAINER_COUNT_MIN (0x00000100)
value TXFS_RM_FLAG_PREFER_AVAILABILITY (0x00020000)
value TXFS_RM_FLAG_PREFER_CONSISTENCY (0x00010000)
value TXFS_RM_FLAG_PRESERVE_CHANGES (0x00002000)
value TXFS_RM_FLAG_RENAME_RM (0x00000002)
value TXFS_RM_FLAG_RESET_RM_AT_NEXT_START (0x00004000)
value TXFS_RM_FLAG_SHRINK_LOG (0x00000800)
value TXFS_RM_STATE_ACTIVE (2)
value TXFS_RM_STATE_NOT_STARTED (0)
value TXFS_RM_STATE_SHUTTING_DOWN (3)
value TXFS_RM_STATE_STARTING (1)
value TXFS_ROLLFORWARD_REDO_FLAG_USE_LAST_REDO_LSN (0x01)
value TXFS_ROLLFORWARD_REDO_FLAG_USE_LAST_VIRTUAL_CLOCK (0x02)
value TXFS_ROLLFORWARD_REDO_VALID_FLAGS ((TXFS_ROLLFORWARD_REDO_FLAG_USE_LAST_REDO_LSN | TXFS_ROLLFORWARD_REDO_FLAG_USE_LAST_VIRTUAL_CLOCK))
value TXFS_SAVEPOINT_CLEAR (0x00000004)
value TXFS_SAVEPOINT_CLEAR_ALL (0x00000010)
value TXFS_SAVEPOINT_ROLLBACK (0x00000002)
value TXFS_SAVEPOINT_SET (0x00000001)
value TXFS_START_RM_FLAG_LOGGING_MODE (0x00000400)
value TXFS_START_RM_FLAG_LOG_AUTO_SHRINK_PERCENTAGE (0x00000020)
value TXFS_START_RM_FLAG_LOG_CONTAINER_COUNT_MAX (0x00000001)
value TXFS_START_RM_FLAG_LOG_CONTAINER_COUNT_MIN (0x00000002)
value TXFS_START_RM_FLAG_LOG_CONTAINER_SIZE (0x00000004)
value TXFS_START_RM_FLAG_LOG_GROWTH_INCREMENT_NUM_CONTAINERS (0x00000008)
value TXFS_START_RM_FLAG_LOG_GROWTH_INCREMENT_PERCENT (0x00000010)
value TXFS_START_RM_FLAG_LOG_NO_CONTAINER_COUNT_MAX (0x00000040)
value TXFS_START_RM_FLAG_LOG_NO_CONTAINER_COUNT_MIN (0x00000080)
value TXFS_START_RM_FLAG_PREFER_AVAILABILITY (0x00002000)
value TXFS_START_RM_FLAG_PREFER_CONSISTENCY (0x00001000)
value TXFS_START_RM_FLAG_PRESERVE_CHANGES (0x00000800)
value TXFS_START_RM_FLAG_RECOVER_BEST_EFFORT (0x00000200)
value TXFS_START_RM_VALID_FLAGS ((TXFS_START_RM_FLAG_LOG_CONTAINER_COUNT_MAX | TXFS_START_RM_FLAG_LOG_CONTAINER_COUNT_MIN | TXFS_START_RM_FLAG_LOG_CONTAINER_SIZE | TXFS_START_RM_FLAG_LOG_GROWTH_INCREMENT_NUM_CONTAINERS | TXFS_START_RM_FLAG_LOG_GROWTH_INCREMENT_PERCENT | TXFS_START_RM_FLAG_LOG_AUTO_SHRINK_PERCENTAGE | TXFS_START_RM_FLAG_RECOVER_BEST_EFFORT | TXFS_START_RM_FLAG_LOG_NO_CONTAINER_COUNT_MAX | TXFS_START_RM_FLAG_LOGGING_MODE | TXFS_START_RM_FLAG_PRESERVE_CHANGES | TXFS_START_RM_FLAG_PREFER_CONSISTENCY | TXFS_START_RM_FLAG_PREFER_AVAILABILITY))
value TXFS_TRANSACTED_VERSION_NONTRANSACTED (0xFFFFFFFE)
value TXFS_TRANSACTED_VERSION_UNCOMMITTED (0xFFFFFFFF)
value TXFS_TRANSACTION_STATE_ACTIVE (0x01)
value TXFS_TRANSACTION_STATE_NONE (0x00)
value TXFS_TRANSACTION_STATE_NOTACTIVE (0x03)
value TXFS_TRANSACTION_STATE_PREPARED (0x02)
value TYPE_E_AMBIGUOUSNAME (_HRESULT_TYPEDEF_(0x8002802CL))
value TYPE_E_BADMODULEKIND (_HRESULT_TYPEDEF_(0x800288BDL))
value TYPE_E_BUFFERTOOSMALL (_HRESULT_TYPEDEF_(0x80028016L))
value TYPE_E_CANTCREATETMPFILE (_HRESULT_TYPEDEF_(0x80028CA3L))
value TYPE_E_CANTLOADLIBRARY (_HRESULT_TYPEDEF_(0x80029C4AL))
value TYPE_E_CIRCULARTYPE (_HRESULT_TYPEDEF_(0x80029C84L))
value TYPE_E_DLLFUNCTIONNOTFOUND (_HRESULT_TYPEDEF_(0x8002802FL))
value TYPE_E_DUPLICATEID (_HRESULT_TYPEDEF_(0x800288C6L))
value TYPE_E_ELEMENTNOTFOUND (_HRESULT_TYPEDEF_(0x8002802BL))
value TYPE_E_FIELDNOTFOUND (_HRESULT_TYPEDEF_(0x80028017L))
value TYPE_E_INCONSISTENTPROPFUNCS (_HRESULT_TYPEDEF_(0x80029C83L))
value TYPE_E_INVALIDID (_HRESULT_TYPEDEF_(0x800288CFL))
value TYPE_E_INVALIDSTATE (_HRESULT_TYPEDEF_(0x80028029L))
value TYPE_E_INVDATAREAD (_HRESULT_TYPEDEF_(0x80028018L))
value TYPE_E_IOERROR (_HRESULT_TYPEDEF_(0x80028CA2L))
value TYPE_E_LIBNOTREGISTERED (_HRESULT_TYPEDEF_(0x8002801DL))
value TYPE_E_NAMECONFLICT (_HRESULT_TYPEDEF_(0x8002802DL))
value TYPE_E_OUTOFBOUNDS (_HRESULT_TYPEDEF_(0x80028CA1L))
value TYPE_E_QUALIFIEDNAMEDISALLOWED (_HRESULT_TYPEDEF_(0x80028028L))
value TYPE_E_REGISTRYACCESS (_HRESULT_TYPEDEF_(0x8002801CL))
value TYPE_E_SIZETOOBIG (_HRESULT_TYPEDEF_(0x800288C5L))
value TYPE_E_TYPEMISMATCH (_HRESULT_TYPEDEF_(0x80028CA0L))
value TYPE_E_UNDEFINEDTYPE (_HRESULT_TYPEDEF_(0x80028027L))
value TYPE_E_UNKNOWNLCID (_HRESULT_TYPEDEF_(0x8002802EL))
value TYPE_E_UNSUPFORMAT (_HRESULT_TYPEDEF_(0x80028019L))
value TYPE_E_WRONGTYPEKIND (_HRESULT_TYPEDEF_(0x8002802AL))
value UAS_EXACTLEGACY (0x00001000)
value UCEERR_BLOCKSFULL (_HRESULT_TYPEDEF_(0x88980409L))
value UCEERR_CHANNELSYNCABANDONED (_HRESULT_TYPEDEF_(0x88980414L))
value UCEERR_CHANNELSYNCTIMEDOUT (_HRESULT_TYPEDEF_(0x88980413L))
value UCEERR_COMMANDTRANSPORTDENIED (_HRESULT_TYPEDEF_(0x88980418L))
value UCEERR_CONNECTIONIDLOOKUPFAILED (_HRESULT_TYPEDEF_(0x88980408L))
value UCEERR_CTXSTACKFRSTTARGETNULL (_HRESULT_TYPEDEF_(0x88980407L))
value UCEERR_FEEDBACK_UNSUPPORTED (_HRESULT_TYPEDEF_(0x88980417L))
value UCEERR_GRAPHICSSTREAMALREADYOPEN (_HRESULT_TYPEDEF_(0x88980420L))
value UCEERR_GRAPHICSSTREAMUNAVAILABLE (_HRESULT_TYPEDEF_(0x88980419L))
value UCEERR_HANDLELOOKUPFAILED (_HRESULT_TYPEDEF_(0x88980405L))
value UCEERR_ILLEGALHANDLE (_HRESULT_TYPEDEF_(0x88980404L))
value UCEERR_ILLEGALPACKET (_HRESULT_TYPEDEF_(0x88980402L))
value UCEERR_ILLEGALRECORDTYPE (_HRESULT_TYPEDEF_(0x8898040CL))
value UCEERR_INVALIDPACKETHEADER (_HRESULT_TYPEDEF_(0x88980400L))
value UCEERR_MALFORMEDPACKET (_HRESULT_TYPEDEF_(0x88980403L))
value UCEERR_MEMORYFAILURE (_HRESULT_TYPEDEF_(0x8898040AL))
value UCEERR_MISSINGBEGINCOMMAND (_HRESULT_TYPEDEF_(0x88980412L))
value UCEERR_MISSINGENDCOMMAND (_HRESULT_TYPEDEF_(0x88980411L))
value UCEERR_NO_MULTIPLE_WORKER_THREADS (_HRESULT_TYPEDEF_(0x8898040FL))
value UCEERR_OUTOFHANDLES (_HRESULT_TYPEDEF_(0x8898040DL))
value UCEERR_PACKETRECORDOUTOFRANGE (_HRESULT_TYPEDEF_(0x8898040BL))
value UCEERR_PARTITION_ZOMBIED (_HRESULT_TYPEDEF_(0x88980423L))
value UCEERR_REMOTINGNOTSUPPORTED (_HRESULT_TYPEDEF_(0x88980410L))
value UCEERR_RENDERTHREADFAILURE (_HRESULT_TYPEDEF_(0x88980406L))
value UCEERR_TRANSPORTDISCONNECTED (_HRESULT_TYPEDEF_(0x88980421L))
value UCEERR_TRANSPORTOVERLOADED (_HRESULT_TYPEDEF_(0x88980422L))
value UCEERR_TRANSPORTUNAVAILABLE (_HRESULT_TYPEDEF_(0x88980416L))
value UCEERR_UNCHANGABLE_UPDATE_ATTEMPTED (_HRESULT_TYPEDEF_(0x8898040EL))
value UCEERR_UNKNOWNPACKET (_HRESULT_TYPEDEF_(0x88980401L))
value UCEERR_UNSUPPORTEDTRANSPORTVERSION (_HRESULT_TYPEDEF_(0x88980415L))
value UCHAR_MAX (0xff)
value UCLEANUI ((SHTDN_REASON_FLAG_CLEAN_UI))
value UDIRTYUI ((SHTDN_REASON_FLAG_DIRTY_UI))
value UILANGUAGE_ENUMPROC (UILANGUAGE_ENUMPROCA)
value UINT_MAX (0xffffffff)
value UISF_ACTIVE (0x4)
value UISF_HIDEACCEL (0x2)
value UISF_HIDEFOCUS (0x1)
value UIS_CLEAR (2)
value UIS_INITIALIZE (3)
value UIS_SET (1)
value UI_CAP_ROTANY (0x00000004)
value UI_E_AMBIGUOUS_MATCH (_HRESULT_TYPEDEF_(0x802A000AL))
value UI_E_BOOLEAN_EXPECTED (_HRESULT_TYPEDEF_(0x802A0008L))
value UI_E_CREATE_FAILED (_HRESULT_TYPEDEF_(0x802A0001L))
value UI_E_DIFFERENT_OWNER (_HRESULT_TYPEDEF_(0x802A0009L))
value UI_E_END_KEYFRAME_NOT_DETERMINED (_HRESULT_TYPEDEF_(0x802A0104L))
value UI_E_FP_OVERFLOW (_HRESULT_TYPEDEF_(0x802A000BL))
value UI_E_ILLEGAL_REENTRANCY (_HRESULT_TYPEDEF_(0x802A0003L))
value UI_E_INVALID_DIMENSION (_HRESULT_TYPEDEF_(0x802A010BL))
value UI_E_INVALID_OUTPUT (_HRESULT_TYPEDEF_(0x802A0007L))
value UI_E_LOOPS_OVERLAP (_HRESULT_TYPEDEF_(0x802A0105L))
value UI_E_OBJECT_SEALED (_HRESULT_TYPEDEF_(0x802A0004L))
value UI_E_PRIMITIVE_OUT_OF_BOUNDS (_HRESULT_TYPEDEF_(0x802A010CL))
value UI_E_SHUTDOWN_CALLED (_HRESULT_TYPEDEF_(0x802A0002L))
value UI_E_START_KEYFRAME_AFTER_END (_HRESULT_TYPEDEF_(0x802A0103L))
value UI_E_STORYBOARD_ACTIVE (_HRESULT_TYPEDEF_(0x802A0101L))
value UI_E_STORYBOARD_NOT_PLAYING (_HRESULT_TYPEDEF_(0x802A0102L))
value UI_E_TIMER_CLIENT_ALREADY_CONNECTED (_HRESULT_TYPEDEF_(0x802A010AL))
value UI_E_TIME_BEFORE_LAST_UPDATE (_HRESULT_TYPEDEF_(0x802A0109L))
value UI_E_TRANSITION_ALREADY_USED (_HRESULT_TYPEDEF_(0x802A0106L))
value UI_E_TRANSITION_ECLIPSED (_HRESULT_TYPEDEF_(0x802A0108L))
value UI_E_TRANSITION_NOT_IN_STORYBOARD (_HRESULT_TYPEDEF_(0x802A0107L))
value UI_E_VALUE_NOT_DETERMINED (_HRESULT_TYPEDEF_(0x802A0006L))
value UI_E_VALUE_NOT_SET (_HRESULT_TYPEDEF_(0x802A0005L))
value UI_E_WINDOW_CLOSED (_HRESULT_TYPEDEF_(0x802A0201L))
value UI_E_WRONG_THREAD (_HRESULT_TYPEDEF_(0x802A000CL))
value ULW_ALPHA (0x00000002)
value ULW_COLORKEY (0x00000001)
value ULW_EX_NORESIZE (0x00000008)
value ULW_OPAQUE (0x00000004)
value UMS_VERSION (RTL_UMS_VERSION)
value UNDEFINE_ALTERNATE (0xD)
value UNDEFINE_PRIMARY (0xC)
value UNICODE_NOCHAR (0xFFFF)
value UNICODE_NULL (((WCHAR)0))
value UNICODE_STRING_MAX_BYTES (((WORD ) 65534))
value UNICODE_STRING_MAX_CHARS ((32767))
value UNIFIEDBUILDREVISION_MIN (0x00000000)
value UNIQUE_NAME (0x00)
value UNIVERSAL_NAME_INFO_LEVEL (0x00000001)
value UNLOAD_DLL_DEBUG_EVENT (7)
value UNLOCK_ELEMENT (1)
value UNPROTECTED_DACL_SECURITY_INFORMATION ((0x20000000L))
value UNPROTECTED_SACL_SECURITY_INFORMATION ((0x10000000L))
value UNRECOVERED_READS_VALID (0x00000008)
value UNRECOVERED_WRITES_VALID (0x00000002)
value UNWIND_CHAIN_LIMIT (32)
value UNWIND_HISTORY_TABLE_SIZE (12)
value UNW_FLAG_CHAININFO (0x4)
value UNW_FLAG_EHANDLER (0x1)
value UNW_FLAG_NHANDLER (0x0)
value UNW_FLAG_NO_EPILOGUE (0x80000000UL)
value UNW_FLAG_UHANDLER (0x2)
value UOI_FLAGS (1)
value UOI_HEAPSIZE (5)
value UOI_IO (6)
value UOI_NAME (2)
value UOI_TIMERPROC_EXCEPTION_SUPPRESSION (7)
value UOI_TYPE (3)
value UOI_USER_SID (4)
value UPDFCACHE_IFBLANK (( 0x10 ))
value UPDFCACHE_IFBLANKORONSAVECACHE (( ( UPDFCACHE_IFBLANK | UPDFCACHE_ONSAVECACHE ) ))
value UPDFCACHE_NODATACACHE (( 0x1 ))
value UPDFCACHE_NORMALCACHE (( 0x8 ))
value UPDFCACHE_ONLYIFBLANK (( 0x80000000 ))
value UPDFCACHE_ONSAVECACHE (( 0x2 ))
value UPDFCACHE_ONSTOPCACHE (( 0x4 ))
value UPDP_CHECK_DRIVERSTORE (0x00000004)
value UPDP_SILENT_UPLOAD (0x00000001)
value UPDP_UPLOAD_ALWAYS (0x00000002)
value URLACTION_ACTIVEX_ALLOW_TDC (0x0000120C)
value URLACTION_ACTIVEX_CONFIRM_NOOBJECTSAFETY (0x00001204)
value URLACTION_ACTIVEX_CURR_MAX (0x0000120C)
value URLACTION_ACTIVEX_DYNSRC_VIDEO_AND_ANIMATION (0x0000120A)
value URLACTION_ACTIVEX_MAX (0x000013ff)
value URLACTION_ACTIVEX_MIN (0x00001200)
value URLACTION_ACTIVEX_NO_WEBOC_SCRIPT (0x00001206)
value URLACTION_ACTIVEX_OVERRIDE_DATA_SAFETY (0x00001202)
value URLACTION_ACTIVEX_OVERRIDE_DOMAINLIST (0x0000120B)
value URLACTION_ACTIVEX_OVERRIDE_OBJECT_SAFETY (0x00001201)
value URLACTION_ACTIVEX_OVERRIDE_OPTIN (0x00001208)
value URLACTION_ACTIVEX_OVERRIDE_REPURPOSEDETECTION (0x00001207)
value URLACTION_ACTIVEX_OVERRIDE_SCRIPT_SAFETY (0x00001203)
value URLACTION_ACTIVEX_RUN (0x00001200)
value URLACTION_ACTIVEX_SCRIPTLET_RUN (0x00001209)
value URLACTION_ACTIVEX_TREATASUNTRUSTED (0x00001205)
value URLACTION_ALLOW_ACTIVEX_FILTERING (0x00002702)
value URLACTION_ALLOW_ANTIMALWARE_SCANNING_OF_ACTIVEX (0x0000270C)
value URLACTION_ALLOW_APEVALUATION (0x00002301)
value URLACTION_ALLOW_AUDIO_VIDEO (0x00002701)
value URLACTION_ALLOW_AUDIO_VIDEO_PLUGINS (0x00002704)
value URLACTION_ALLOW_CROSSDOMAIN_APPCACHE_MANIFEST (0x0000270A)
value URLACTION_ALLOW_CROSSDOMAIN_DROP_ACROSS_WINDOWS (0x00002709)
value URLACTION_ALLOW_CROSSDOMAIN_DROP_WITHIN_WINDOW (0x00002708)
value URLACTION_ALLOW_CSS_EXPRESSIONS (0x0000270D)
value URLACTION_ALLOW_JSCRIPT_IE (0x0000140D)
value URLACTION_ALLOW_RENDER_LEGACY_DXTFILTERS (0x0000270B)
value URLACTION_ALLOW_RESTRICTEDPROTOCOLS (0x00002300)
value URLACTION_ALLOW_STRUCTURED_STORAGE_SNIFFING (0x00002703)
value URLACTION_ALLOW_VBSCRIPT_IE (0x0000140C)
value URLACTION_ALLOW_XDOMAIN_SUBFRAME_RESIZE (0x00001408)
value URLACTION_ALLOW_XHR_EVALUATION (0x00002302)
value URLACTION_ALLOW_ZONE_ELEVATION_OPT_OUT_ADDITION (0x00002706)
value URLACTION_ALLOW_ZONE_ELEVATION_VIA_OPT_OUT (0x00002705)
value URLACTION_AUTHENTICATE_CLIENT (0x00001A01)
value URLACTION_AUTOMATIC_ACTIVEX_UI (0x00002201)
value URLACTION_AUTOMATIC_DOWNLOAD_UI (0x00002200)
value URLACTION_AUTOMATIC_DOWNLOAD_UI_MIN (0x00002200)
value URLACTION_BEHAVIOR_MIN (0x00002000)
value URLACTION_BEHAVIOR_RUN (0x00002000)
value URLACTION_CHANNEL_SOFTDIST_MAX (0x00001Eff)
value URLACTION_CHANNEL_SOFTDIST_MIN (0x00001E00)
value URLACTION_CHANNEL_SOFTDIST_PERMISSIONS (0x00001E05)
value URLACTION_CLIENT_CERT_PROMPT (0x00001A04)
value URLACTION_COOKIES (0x00001A02)
value URLACTION_COOKIES_ENABLED (0x00001A10)
value URLACTION_COOKIES_SESSION (0x00001A03)
value URLACTION_COOKIES_SESSION_THIRD_PARTY (0x00001A06)
value URLACTION_COOKIES_THIRD_PARTY (0x00001A05)
value URLACTION_CREDENTIALS_USE (0x00001A00)
value URLACTION_CROSS_DOMAIN_DATA (0x00001406)
value URLACTION_DOTNET_USERCONTROLS (0x00002005)
value URLACTION_DOWNLOAD_CURR_MAX (0x00001004)
value URLACTION_DOWNLOAD_MAX (0x000011FF)
value URLACTION_DOWNLOAD_MIN (0x00001000)
value URLACTION_DOWNLOAD_SIGNED_ACTIVEX (0x00001001)
value URLACTION_DOWNLOAD_UNSIGNED_ACTIVEX (0x00001004)
value URLACTION_FEATURE_BLOCK_INPUT_PROMPTS (0x00002105)
value URLACTION_FEATURE_CROSSDOMAIN_FOCUS_CHANGE (0x00002107)
value URLACTION_FEATURE_DATA_BINDING (0x00002106)
value URLACTION_FEATURE_FORCE_ADDR_AND_STATUS (0x00002104)
value URLACTION_FEATURE_MIME_SNIFFING (0x00002100)
value URLACTION_FEATURE_MIN (0x00002100)
value URLACTION_FEATURE_SCRIPT_STATUS_BAR (0x00002103)
value URLACTION_FEATURE_WINDOW_RESTRICTIONS (0x00002102)
value URLACTION_FEATURE_ZONE_ELEVATION (0x00002101)
value URLACTION_HTML_ALLOW_CROSS_DOMAIN_CANVAS (0x0000160D)
value URLACTION_HTML_ALLOW_CROSS_DOMAIN_TEXTTRACK (0x00001610)
value URLACTION_HTML_ALLOW_CROSS_DOMAIN_WEBWORKER (0x0000160F)
value URLACTION_HTML_ALLOW_INDEXEDDB (0x00001611)
value URLACTION_HTML_ALLOW_INJECTED_DYNAMIC_HTML (0x0000160B)
value URLACTION_HTML_ALLOW_WINDOW_CLOSE (0x0000160E)
value URLACTION_HTML_FONT_DOWNLOAD (0x00001604)
value URLACTION_HTML_INCLUDE_FILE_PATH (0x0000160A)
value URLACTION_HTML_JAVA_RUN (0x00001605)
value URLACTION_HTML_MAX (0x000017ff)
value URLACTION_HTML_META_REFRESH (0x00001608)
value URLACTION_HTML_MIN (0x00001600)
value URLACTION_HTML_MIXED_CONTENT (0x00001609)
value URLACTION_HTML_SUBFRAME_NAVIGATE (0x00001607)
value URLACTION_HTML_SUBMIT_FORMS (0x00001601)
value URLACTION_HTML_SUBMIT_FORMS_FROM (0x00001602)
value URLACTION_HTML_SUBMIT_FORMS_TO (0x00001603)
value URLACTION_HTML_USERDATA_SAVE (0x00001606)
value URLACTION_INFODELIVERY_CURR_MAX (0x00001D06)
value URLACTION_INFODELIVERY_MAX (0x00001Dff)
value URLACTION_INFODELIVERY_MIN (0x00001D00)
value URLACTION_INFODELIVERY_NO_ADDING_CHANNELS (0x00001D00)
value URLACTION_INFODELIVERY_NO_ADDING_SUBSCRIPTIONS (0x00001D03)
value URLACTION_INFODELIVERY_NO_CHANNEL_LOGGING (0x00001D06)
value URLACTION_INFODELIVERY_NO_EDITING_CHANNELS (0x00001D01)
value URLACTION_INFODELIVERY_NO_EDITING_SUBSCRIPTIONS (0x00001D04)
value URLACTION_INFODELIVERY_NO_REMOVING_CHANNELS (0x00001D02)
value URLACTION_INFODELIVERY_NO_REMOVING_SUBSCRIPTIONS (0x00001D05)
value URLACTION_INPRIVATE_BLOCKING (0x00002700)
value URLACTION_JAVA_CURR_MAX (0x00001C00)
value URLACTION_JAVA_MAX (0x00001Cff)
value URLACTION_JAVA_MIN (0x00001C00)
value URLACTION_JAVA_PERMISSIONS (0x00001C00)
value URLACTION_LOOSE_XAML (0x00002402)
value URLACTION_LOWRIGHTS (0x00002500)
value URLACTION_MIN (0x00001000)
value URLACTION_NETWORK_CURR_MAX (0x00001A10)
value URLACTION_NETWORK_MAX (0x00001Bff)
value URLACTION_NETWORK_MIN (0x00001A00)
value URLACTION_PLUGGABLE_PROTOCOL_XHR (0x0000140B)
value URLACTION_SCRIPT_CURR_MAX (0x0000140D)
value URLACTION_SCRIPT_JAVA_USE (0x00001402)
value URLACTION_SCRIPT_MAX (0x000015ff)
value URLACTION_SCRIPT_MIN (0x00001400)
value URLACTION_SCRIPT_NAVIGATE (0x0000140A)
value URLACTION_SCRIPT_OVERRIDE_SAFETY (0x00001401)
value URLACTION_SCRIPT_PASTE (0x00001407)
value URLACTION_SCRIPT_RUN (0x00001400)
value URLACTION_SCRIPT_SAFE_ACTIVEX (0x00001405)
value URLACTION_SCRIPT_XSSFILTER (0x00001409)
value URLACTION_SHELL_ALLOW_CROSS_SITE_SHARE (0x00001811)
value URLACTION_SHELL_CURR_MAX (0x00001812)
value URLACTION_SHELL_ENHANCED_DRAGDROP_SECURITY (0x0000180B)
value URLACTION_SHELL_EXECUTE_HIGHRISK (0x00001806)
value URLACTION_SHELL_EXECUTE_LOWRISK (0x00001808)
value URLACTION_SHELL_EXECUTE_MODRISK (0x00001807)
value URLACTION_SHELL_EXTENSIONSECURITY (0x0000180C)
value URLACTION_SHELL_FILE_DOWNLOAD (0x00001803)
value URLACTION_SHELL_INSTALL_DTITEMS (0x00001800)
value URLACTION_SHELL_MAX (0x000019ff)
value URLACTION_SHELL_MIN (0x00001800)
value URLACTION_SHELL_MOVE_OR_COPY (0x00001802)
value URLACTION_SHELL_POPUPMGR (0x00001809)
value URLACTION_SHELL_PREVIEW (0x0000180F)
value URLACTION_SHELL_REMOTEQUERY (0x0000180E)
value URLACTION_SHELL_RTF_OBJECTS_LOAD (0x0000180A)
value URLACTION_SHELL_SECURE_DRAGSOURCE (0x0000180D)
value URLACTION_SHELL_SHARE (0x00001810)
value URLACTION_SHELL_SHELLEXECUTE (0x00001806)
value URLACTION_SHELL_TOCTOU_RISK (0x00001812)
value URLACTION_SHELL_VERB (0x00001804)
value URLACTION_SHELL_WEBVIEW_VERB (0x00001805)
value URLACTION_WINDOWS_BROWSER_APPLICATIONS (0x00002400)
value URLACTION_WINFX_SETUP (0x00002600)
value URLACTION_XPS_DOCUMENTS (0x00002401)
value URLMON_OPTION_URL_ENCODING (0x10000004)
value URLMON_OPTION_USERAGENT (0x10000001)
value URLMON_OPTION_USERAGENT_REFRESH (0x10000002)
value URLMON_OPTION_USE_BINDSTRINGCREDS (0x10000008)
value URLMON_OPTION_USE_BROWSERAPPSDOCUMENTS (0x10000010)
value URLOSTRM_GETNEWESTVERSION (0x3)
value URLOSTRM_USECACHEDCOPY (0x2)
value URLOSTRM_USECACHEDCOPY_ONLY (0x1)
value URLPOLICY_ACTIVEX_CHECK_LIST (0x00010000)
value URLPOLICY_ALLOW (0x00)
value URLPOLICY_AUTHENTICATE_CHALLENGE_RESPONSE (0x00010000)
value URLPOLICY_AUTHENTICATE_CLEARTEXT_OK (0x00000000)
value URLPOLICY_AUTHENTICATE_MUTUAL_ONLY (0x00030000)
value URLPOLICY_BEHAVIOR_CHECK_LIST (0x00010000)
value URLPOLICY_CHANNEL_SOFTDIST_AUTOINSTALL (0x00030000)
value URLPOLICY_CHANNEL_SOFTDIST_PRECACHE (0x00020000)
value URLPOLICY_CHANNEL_SOFTDIST_PROHIBIT (0x00010000)
value URLPOLICY_CREDENTIALS_ANONYMOUS_ONLY (0x00030000)
value URLPOLICY_CREDENTIALS_CONDITIONAL_PROMPT (0x00020000)
value URLPOLICY_CREDENTIALS_MUST_PROMPT_USER (0x00010000)
value URLPOLICY_CREDENTIALS_SILENT_LOGON_OK (0x00000000)
value URLPOLICY_DISALLOW (0x03)
value URLPOLICY_DONTCHECKDLGBOX (0x100)
value URLPOLICY_JAVA_CUSTOM (0x00800000)
value URLPOLICY_JAVA_HIGH (0x00010000)
value URLPOLICY_JAVA_LOW (0x00030000)
value URLPOLICY_JAVA_MEDIUM (0x00020000)
value URLPOLICY_JAVA_PROHIBIT (0x00000000)
value URLPOLICY_LOG_ON_ALLOW (0x40)
value URLPOLICY_LOG_ON_DISALLOW (0x80)
value URLPOLICY_MASK_PERMISSIONS (0x0f)
value URLPOLICY_NOTIFY_ON_ALLOW (0x10)
value URLPOLICY_NOTIFY_ON_DISALLOW (0x20)
value URLPOLICY_QUERY (0x01)
value URLZONE_ESC_FLAG (0x100)
value URL_MK_LEGACY (0)
value URL_MK_NO_CANONICALIZE (2)
value URL_MK_UNIFORM (1)
value URL_OID_CERTIFICATE_CRL_DIST_POINT (((LPCSTR)2))
value URL_OID_CERTIFICATE_CRL_DIST_POINT_AND_OCSP (((LPCSTR)11))
value URL_OID_CERTIFICATE_FRESHEST_CRL (((LPCSTR)6))
value URL_OID_CERTIFICATE_ISSUER (((LPCSTR)1))
value URL_OID_CERTIFICATE_OCSP (((LPCSTR)9))
value URL_OID_CERTIFICATE_OCSP_AND_CRL_DIST_POINT (((LPCSTR)10))
value URL_OID_CERTIFICATE_ONLY_OCSP (((LPCSTR)13))
value URL_OID_CRL_FRESHEST_CRL (((LPCSTR)7))
value URL_OID_CRL_ISSUER (((LPCSTR)5))
value URL_OID_CROSS_CERT_DIST_POINT (((LPCSTR)8))
value URL_OID_CROSS_CERT_SUBJECT_INFO_ACCESS (((LPCSTR)12))
value URL_OID_CTL_ISSUER (((LPCSTR)3))
value URL_OID_CTL_NEXT_UPDATE (((LPCSTR)4))
value USAGE_MATCH_TYPE_AND (0x00000000)
value USAGE_MATCH_TYPE_OR (0x00000001)
value USER_CALL_IS_ASYNC (0x0100)
value USER_CALL_NEW_CORRELATION_DESC (0x0200)
value USER_CET_ENVIRONMENT_VBS_BASIC_ENCLAVE (0x00000011)
value USER_CET_ENVIRONMENT_VBS_ENCLAVE (0x00000010)
value USER_DEFAULT_SCREEN_DPI (96)
value USER_MARSHAL_FC_BYTE (1)
value USER_MARSHAL_FC_CHAR (2)
value USER_MARSHAL_FC_DOUBLE (12)
value USER_MARSHAL_FC_FLOAT (10)
value USER_MARSHAL_FC_HYPER (11)
value USER_MARSHAL_FC_LONG (8)
value USER_MARSHAL_FC_SHORT (6)
value USER_MARSHAL_FC_SMALL (3)
value USER_MARSHAL_FC_ULONG (9)
value USER_MARSHAL_FC_USHORT (7)
value USER_MARSHAL_FC_USMALL (4)
value USER_MARSHAL_FC_WCHAR (5)
value USER_TIMER_MAXIMUM (0x7FFFFFFF)
value USER_TIMER_MINIMUM (0x0000000A)
value USHRT_MAX (0xffff)
value USN_DELETE_FLAG_DELETE ((0x00000001))
value USN_DELETE_FLAG_NOTIFY ((0x00000002))
value USN_DELETE_VALID_FLAGS ((0x00000003))
value USN_PAGE_SIZE ((0x1000))
value USN_REASON_BASIC_INFO_CHANGE ((0x00008000))
value USN_REASON_CLOSE ((0x80000000))
value USN_REASON_COMPRESSION_CHANGE ((0x00020000))
value USN_REASON_DATA_EXTEND ((0x00000002))
value USN_REASON_DATA_OVERWRITE ((0x00000001))
value USN_REASON_DATA_TRUNCATION ((0x00000004))
value USN_REASON_DESIRED_STORAGE_CLASS_CHANGE ((0x01000000))
value USN_REASON_EA_CHANGE ((0x00000400))
value USN_REASON_ENCRYPTION_CHANGE ((0x00040000))
value USN_REASON_FILE_CREATE ((0x00000100))
value USN_REASON_FILE_DELETE ((0x00000200))
value USN_REASON_HARD_LINK_CHANGE ((0x00010000))
value USN_REASON_INDEXABLE_CHANGE ((0x00004000))
value USN_REASON_INTEGRITY_CHANGE ((0x00800000))
value USN_REASON_NAMED_DATA_EXTEND ((0x00000020))
value USN_REASON_NAMED_DATA_OVERWRITE ((0x00000010))
value USN_REASON_NAMED_DATA_TRUNCATION ((0x00000040))
value USN_REASON_OBJECT_ID_CHANGE ((0x00080000))
value USN_REASON_RENAME_NEW_NAME ((0x00002000))
value USN_REASON_RENAME_OLD_NAME ((0x00001000))
value USN_REASON_REPARSE_POINT_CHANGE ((0x00100000))
value USN_REASON_SECURITY_CHANGE ((0x00000800))
value USN_REASON_STREAM_CHANGE ((0x00200000))
value USN_REASON_TRANSACTED_CHANGE ((0x00400000))
value USN_SOURCE_AUXILIARY_DATA ((0x00000002))
value USN_SOURCE_CLIENT_REPLICATION_MANAGEMENT ((0x00000008))
value USN_SOURCE_DATA_MANAGEMENT ((0x00000001))
value USN_SOURCE_REPLICATION_MANAGEMENT ((0x00000004))
value USN_SOURCE_VALID_FLAGS ((USN_SOURCE_DATA_MANAGEMENT | USN_SOURCE_AUXILIARY_DATA | USN_SOURCE_REPLICATION_MANAGEMENT | USN_SOURCE_CLIENT_REPLICATION_MANAGEMENT))
value UTC_E_ACTION_NOT_SUPPORTED_IN_DESTINATION (_HRESULT_TYPEDEF_(0x87C51044L))
value UTC_E_AGENT_DIAGNOSTICS_TOO_LARGE (_HRESULT_TYPEDEF_(0x87C51055L))
value UTC_E_ALTERNATIVE_TRACE_CANNOT_PREEMPT (_HRESULT_TYPEDEF_(0x87C51002L))
value UTC_E_AOT_NOT_RUNNING (_HRESULT_TYPEDEF_(0x87C51003L))
value UTC_E_API_BUSY (_HRESULT_TYPEDEF_(0x87C5102BL))
value UTC_E_API_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x87C5103CL))
value UTC_E_API_RESULT_UNAVAILABLE (_HRESULT_TYPEDEF_(0x87C51028L))
value UTC_E_BINARY_MISSING (_HRESULT_TYPEDEF_(0x87C51034L))
value UTC_E_CANNOT_LOAD_SCENARIO_EDITOR_XML (_HRESULT_TYPEDEF_(0x87C5101FL))
value UTC_E_CERT_REV_FAILED (_HRESULT_TYPEDEF_(0x87C5103FL))
value UTC_E_CHILD_PROCESS_FAILED (_HRESULT_TYPEDEF_(0x87C5101DL))
value UTC_E_COMMAND_LINE_NOT_AUTHORIZED (_HRESULT_TYPEDEF_(0x87C5101EL))
value UTC_E_DELAY_TERMINATED (_HRESULT_TYPEDEF_(0x87C51025L))
value UTC_E_DEVICE_TICKET_ERROR (_HRESULT_TYPEDEF_(0x87C51026L))
value UTC_E_DIAGRULES_SCHEMAVERSION_MISMATCH (_HRESULT_TYPEDEF_(0x87C5100AL))
value UTC_E_ESCALATION_ALREADY_RUNNING (_HRESULT_TYPEDEF_(0x87C5100FL))
value UTC_E_ESCALATION_CANCELLED_AT_SHUTDOWN (_HRESULT_TYPEDEF_(0x87C5105AL))
value UTC_E_ESCALATION_DIRECTORY_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x87C5102FL))
value UTC_E_ESCALATION_NOT_AUTHORIZED (_HRESULT_TYPEDEF_(0x87C5101BL))
value UTC_E_ESCALATION_TIMED_OUT (_HRESULT_TYPEDEF_(0x87C51020L))
value UTC_E_EVENTLOG_ENTRY_MALFORMED (_HRESULT_TYPEDEF_(0x87C51009L))
value UTC_E_EXCLUSIVITY_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x87C5102DL))
value UTC_E_EXE_TERMINATED (_HRESULT_TYPEDEF_(0x87C5101AL))
value UTC_E_FAILED_TO_RECEIVE_AGENT_DIAGNOSTICS (_HRESULT_TYPEDEF_(0x87C51056L))
value UTC_E_FAILED_TO_RESOLVE_CONTAINER_ID (_HRESULT_TYPEDEF_(0x87C51036L))
value UTC_E_FAILED_TO_START_NDISCAP (_HRESULT_TYPEDEF_(0x87C51040L))
value UTC_E_FILTER_FUNCTION_RESTRICTED (_HRESULT_TYPEDEF_(0x87C51048L))
value UTC_E_FILTER_ILLEGAL_EVAL (_HRESULT_TYPEDEF_(0x87C51053L))
value UTC_E_FILTER_INVALID_COMMAND (_HRESULT_TYPEDEF_(0x87C51052L))
value UTC_E_FILTER_INVALID_FUNCTION (_HRESULT_TYPEDEF_(0x87C51050L))
value UTC_E_FILTER_INVALID_FUNCTION_PARAMS (_HRESULT_TYPEDEF_(0x87C51051L))
value UTC_E_FILTER_INVALID_TYPE (_HRESULT_TYPEDEF_(0x87C51046L))
value UTC_E_FILTER_MISSING_ATTRIBUTE (_HRESULT_TYPEDEF_(0x87C51045L))
value UTC_E_FILTER_VARIABLE_NOT_FOUND (_HRESULT_TYPEDEF_(0x87C51047L))
value UTC_E_FILTER_VERSION_MISMATCH (_HRESULT_TYPEDEF_(0x87C51049L))
value UTC_E_FORWARDER_ALREADY_DISABLED (_HRESULT_TYPEDEF_(0x87C51008L))
value UTC_E_FORWARDER_ALREADY_ENABLED (_HRESULT_TYPEDEF_(0x87C51007L))
value UTC_E_FORWARDER_PRODUCER_MISMATCH (_HRESULT_TYPEDEF_(0x87C51012L))
value UTC_E_GETFILEINFOACTION_FILE_NOT_APPROVED (_HRESULT_TYPEDEF_(0x87C5105BL))
value UTC_E_GETFILE_EXTERNAL_PATH_NOT_APPROVED (_HRESULT_TYPEDEF_(0x87C5103DL))
value UTC_E_GETFILE_FILE_PATH_NOT_APPROVED (_HRESULT_TYPEDEF_(0x87C5102EL))
value UTC_E_INSUFFICIENT_SPACE_TO_START_TRACE (_HRESULT_TYPEDEF_(0x87C51059L))
value UTC_E_INTENTIONAL_SCRIPT_FAILURE (_HRESULT_TYPEDEF_(0x87C51013L))
value UTC_E_INVALID_AGGREGATION_STRUCT (_HRESULT_TYPEDEF_(0x87C51043L))
value UTC_E_INVALID_CUSTOM_FILTER (_HRESULT_TYPEDEF_(0x87C5100CL))
value UTC_E_INVALID_FILTER (_HRESULT_TYPEDEF_(0x87C51019L))
value UTC_E_KERNELDUMP_LIMIT_REACHED (_HRESULT_TYPEDEF_(0x87C51041L))
value UTC_E_MISSING_AGGREGATE_EVENT_TAG (_HRESULT_TYPEDEF_(0x87C51042L))
value UTC_E_MULTIPLE_TIME_TRIGGER_ON_SINGLE_STATE (_HRESULT_TYPEDEF_(0x87C51033L))
value UTC_E_NO_WER_LOGGER_SUPPORTED (_HRESULT_TYPEDEF_(0x87C51015L))
value UTC_E_PERFTRACK_ALREADY_TRACING (_HRESULT_TYPEDEF_(0x87C51010L))
value UTC_E_REACHED_MAX_ESCALATIONS (_HRESULT_TYPEDEF_(0x87C51011L))
value UTC_E_REESCALATED_TOO_QUICKLY (_HRESULT_TYPEDEF_(0x87C5100EL))
value UTC_E_RPC_TIMEOUT (_HRESULT_TYPEDEF_(0x87C51029L))
value UTC_E_RPC_WAIT_FAILED (_HRESULT_TYPEDEF_(0x87C5102AL))
value UTC_E_SCENARIODEF_NOT_FOUND (_HRESULT_TYPEDEF_(0x87C51005L))
value UTC_E_SCENARIODEF_SCHEMAVERSION_MISMATCH (_HRESULT_TYPEDEF_(0x87C51018L))
value UTC_E_SCENARIO_HAS_NO_ACTIONS (_HRESULT_TYPEDEF_(0x87C51057L))
value UTC_E_SCENARIO_THROTTLED (_HRESULT_TYPEDEF_(0x87C5103BL))
value UTC_E_SCRIPT_MISSING (_HRESULT_TYPEDEF_(0x87C5103AL))
value UTC_E_SCRIPT_TERMINATED (_HRESULT_TYPEDEF_(0x87C5100BL))
value UTC_E_SCRIPT_TYPE_INVALID (_HRESULT_TYPEDEF_(0x87C51004L))
value UTC_E_SETREGKEYACTION_TYPE_NOT_APPROVED (_HRESULT_TYPEDEF_(0x87C5105CL))
value UTC_E_SETUP_NOT_AUTHORIZED (_HRESULT_TYPEDEF_(0x87C5101CL))
value UTC_E_SETUP_TIMED_OUT (_HRESULT_TYPEDEF_(0x87C51021L))
value UTC_E_SIF_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x87C51024L))
value UTC_E_SQM_INIT_FAILED (_HRESULT_TYPEDEF_(0x87C51014L))
value UTC_E_THROTTLED (_HRESULT_TYPEDEF_(0x87C51038L))
value UTC_E_TIME_TRIGGER_INVALID_TIME_RANGE (_HRESULT_TYPEDEF_(0x87C51032L))
value UTC_E_TIME_TRIGGER_ONLY_VALID_ON_SINGLE_TRANSITION (_HRESULT_TYPEDEF_(0x87C51031L))
value UTC_E_TIME_TRIGGER_ON_START_INVALID (_HRESULT_TYPEDEF_(0x87C51030L))
value UTC_E_TOGGLE_TRACE_STARTED (_HRESULT_TYPEDEF_(0x87C51001L))
value UTC_E_TRACEPROFILE_NOT_FOUND (_HRESULT_TYPEDEF_(0x87C51006L))
value UTC_E_TRACERS_DONT_EXIST (_HRESULT_TYPEDEF_(0x87C51016L))
value UTC_E_TRACE_BUFFER_LIMIT_EXCEEDED (_HRESULT_TYPEDEF_(0x87C51027L))
value UTC_E_TRACE_MIN_DURATION_REQUIREMENT_NOT_MET (_HRESULT_TYPEDEF_(0x87C5102CL))
value UTC_E_TRACE_NOT_RUNNING (_HRESULT_TYPEDEF_(0x87C5100DL))
value UTC_E_TRACE_THROTTLED (_HRESULT_TYPEDEF_(0x87C5105DL))
value UTC_E_TRIGGER_MISMATCH (_HRESULT_TYPEDEF_(0x87C51022L))
value UTC_E_TRIGGER_NOT_FOUND (_HRESULT_TYPEDEF_(0x87C51023L))
value UTC_E_TRY_GET_SCENARIO_TIMEOUT_EXCEEDED (_HRESULT_TYPEDEF_(0x87C5103EL))
value UTC_E_TTTRACER_RETURNED_ERROR (_HRESULT_TYPEDEF_(0x87C51054L))
value UTC_E_TTTRACER_STORAGE_FULL (_HRESULT_TYPEDEF_(0x87C51058L))
value UTC_E_UNABLE_TO_RESOLVE_SESSION (_HRESULT_TYPEDEF_(0x87C51037L))
value UTC_E_UNAPPROVED_SCRIPT (_HRESULT_TYPEDEF_(0x87C51039L))
value UTC_E_WINRT_INIT_FAILED (_HRESULT_TYPEDEF_(0x87C51017L))
value VALID_INHERIT_FLAGS ((0x1F))
value VALID_NTFT (0xC0)
value VALID_WRITE_USN_REASON_MASK ((USN_REASON_DATA_OVERWRITE | USN_REASON_CLOSE))
value VARCMP_EQ (1)
value VARCMP_GT (2)
value VARCMP_LT (0)
value VARCMP_NULL (3)
value VARIABLE_PITCH (2)
value VARIANT_ALPHABOOL (0x02)
value VARIANT_CALENDAR_GREGORIAN (0x40)
value VARIANT_CALENDAR_HIJRI (0x08)
value VARIANT_CALENDAR_THAI (0x20)
value VARIANT_FALSE (((VARIANT_BOOL)0))
value VARIANT_LOCALBOOL (0x10)
value VARIANT_NOUSEROVERRIDE (0x04)
value VARIANT_NOVALUEPROP (0x01)
value VARIANT_TRUE (((VARIANT_BOOL)-1))
value VARIANT_USE_NLS (0x80)
value VAR_CALENDAR_GREGORIAN (((DWORD)0x00000100))
value VAR_CALENDAR_HIJRI (((DWORD)0x00000008))
value VAR_CALENDAR_THAI (((DWORD)0x00000080))
value VAR_DATEVALUEONLY (((DWORD)0x00000002))
value VAR_FORMAT_NOSUBSTITUTE (((DWORD)0x00000020))
value VAR_FOURDIGITYEARS (((DWORD)0x00000040))
value VAR_LOCALBOOL (((DWORD)0x00000010))
value VAR_TIMEVALUEONLY (((DWORD)0x00000001))
value VAR_VALIDDATE (((DWORD)0x00000004))
value VBS_BASIC_PAGE_MEASURED_DATA (0x00000001)
value VBS_BASIC_PAGE_SYSTEM_CALL (0x00000005)
value VBS_BASIC_PAGE_THREAD_DESCRIPTOR (0x00000004)
value VBS_BASIC_PAGE_UNMEASURED_DATA (0x00000002)
value VBS_BASIC_PAGE_ZERO_FILL (0x00000003)
value VENDOR_ID_LENGTH (8)
value VERTRES (10)
value VERTSIZE (6)
value VER_AND (6)
value VER_BUILDNUMBER (0x0000004)
value VER_CONDITION_MASK (7)
value VER_EQUAL (1)
value VER_GREATER (2)
value VER_GREATER_EQUAL (3)
value VER_LESS (4)
value VER_LESS_EQUAL (5)
value VER_MAJORVERSION (0x0000002)
value VER_MINORVERSION (0x0000001)
value VER_NT_DOMAIN_CONTROLLER (0x0000002)
value VER_NT_SERVER (0x0000003)
value VER_NT_WORKSTATION (0x0000001)
value VER_NUM_BITS_PER_CONDITION_MASK (3)
value VER_OR (7)
value VER_PLATFORMID (0x0000008)
value VER_PRODUCT_TYPE (0x0000080)
value VER_SERVER_NT (0x80000000)
value VER_SERVICEPACKMAJOR (0x0000020)
value VER_SERVICEPACKMINOR (0x0000010)
value VER_SUITENAME (0x0000040)
value VER_SUITE_BACKOFFICE (0x00000004)
value VER_SUITE_BLADE (0x00000400)
value VER_SUITE_COMMUNICATIONS (0x00000008)
value VER_SUITE_COMPUTE_SERVER (0x00004000)
value VER_SUITE_DATACENTER (0x00000080)
value VER_SUITE_EMBEDDEDNT (0x00000040)
value VER_SUITE_EMBEDDED_RESTRICTED (0x00000800)
value VER_SUITE_ENTERPRISE (0x00000002)
value VER_SUITE_MULTIUSERTS (0x00020000)
value VER_SUITE_PERSONAL (0x00000200)
value VER_SUITE_SECURITY_APPLIANCE (0x00001000)
value VER_SUITE_SINGLEUSERTS (0x00000100)
value VER_SUITE_SMALLBUSINESS (0x00000001)
value VER_SUITE_SMALLBUSINESS_RESTRICTED (0x00000020)
value VER_SUITE_STORAGE_SERVER (0x00002000)
value VER_SUITE_TERMINAL (0x00000010)
value VER_SUITE_WH_SERVER (0x00008000)
value VER_WORKSTATION_NT (0x40000000)
value VFFF_ISSHAREDFILE (0x0001)
value VFF_BUFFTOOSMALL (0x0004)
value VFF_CURNEDEST (0x0001)
value VFF_FILEINUSE (0x0002)
value VFT_APP (0x00000001L)
value VFT_DLL (0x00000002L)
value VFT_DRV (0x00000003L)
value VFT_FONT (0x00000004L)
value VFT_STATIC_LIB (0x00000007L)
value VFT_UNKNOWN (0x00000000L)
value VFT_VXD (0x00000005L)
value VIETNAMESE_CHARSET (163)
value VIEW_E_DRAW (_HRESULT_TYPEDEF_(0x80040140L))
value VIEW_E_FIRST (0x80040140L)
value VIEW_E_LAST (0x8004014FL)
value VIEW_S_ALREADY_FROZEN (_HRESULT_TYPEDEF_(0x00040140L))
value VIEW_S_FIRST (0x00040140L)
value VIEW_S_LAST (0x0004014FL)
value VIFF_DONTDELETEOLD (0x0002)
value VIFF_FORCEINSTALL (0x0001)
value VIF_ACCESSVIOLATION (0x00000200L)
value VIF_BUFFTOOSMALL (0x00040000L)
value VIF_CANNOTCREATE (0x00000800L)
value VIF_CANNOTDELETE (0x00001000L)
value VIF_CANNOTDELETECUR (0x00004000L)
value VIF_CANNOTLOADCABINET (0x00100000L)
value VIF_CANNOTREADDST (0x00020000L)
value VIF_CANNOTREADSRC (0x00010000L)
value VIF_CANNOTRENAME (0x00002000L)
value VIF_DIFFCODEPG (0x00000010L)
value VIF_DIFFLANG (0x00000008L)
value VIF_DIFFTYPE (0x00000020L)
value VIF_FILEINUSE (0x00000080L)
value VIF_MISMATCH (0x00000002L)
value VIF_OUTOFMEMORY (0x00008000L)
value VIF_OUTOFSPACE (0x00000100L)
value VIF_SHARINGVIOLATION (0x00000400L)
value VIF_SRCOLD (0x00000004L)
value VIF_TEMPFILE (0x00000001L)
value VIF_WRITEPROT (0x00000040L)
value VK_ACCEPT (0x1E)
value VK_ADD (0x6B)
value VK_APPS (0x5D)
value VK_ATTN (0xF6)
value VK_BACK (0x08)
value VK_BROWSER_BACK (0xA6)
value VK_BROWSER_FAVORITES (0xAB)
value VK_BROWSER_FORWARD (0xA7)
value VK_BROWSER_HOME (0xAC)
value VK_BROWSER_REFRESH (0xA8)
value VK_BROWSER_SEARCH (0xAA)
value VK_BROWSER_STOP (0xA9)
value VK_CANCEL (0x03)
value VK_CAPITAL (0x14)
value VK_CLEAR (0x0C)
value VK_CONTROL (0x11)
value VK_CONVERT (0x1C)
value VK_CRSEL (0xF7)
value VK_DECIMAL (0x6E)
value VK_DELETE (0x2E)
value VK_DIVIDE (0x6F)
value VK_DOWN (0x28)
value VK_END (0x23)
value VK_EREOF (0xF9)
value VK_ESCAPE (0x1B)
value VK_EXECUTE (0x2B)
value VK_EXSEL (0xF8)
value VK_FINAL (0x18)
value VK_GAMEPAD_A (0xC3)
value VK_GAMEPAD_B (0xC4)
value VK_GAMEPAD_DPAD_DOWN (0xCC)
value VK_GAMEPAD_DPAD_LEFT (0xCD)
value VK_GAMEPAD_DPAD_RIGHT (0xCE)
value VK_GAMEPAD_DPAD_UP (0xCB)
value VK_GAMEPAD_LEFT_SHOULDER (0xC8)
value VK_GAMEPAD_LEFT_THUMBSTICK_BUTTON (0xD1)
value VK_GAMEPAD_LEFT_THUMBSTICK_DOWN (0xD4)
value VK_GAMEPAD_LEFT_THUMBSTICK_LEFT (0xD6)
value VK_GAMEPAD_LEFT_THUMBSTICK_RIGHT (0xD5)
value VK_GAMEPAD_LEFT_THUMBSTICK_UP (0xD3)
value VK_GAMEPAD_LEFT_TRIGGER (0xC9)
value VK_GAMEPAD_MENU (0xCF)
value VK_GAMEPAD_RIGHT_SHOULDER (0xC7)
value VK_GAMEPAD_RIGHT_THUMBSTICK_BUTTON (0xD2)
value VK_GAMEPAD_RIGHT_THUMBSTICK_DOWN (0xD8)
value VK_GAMEPAD_RIGHT_THUMBSTICK_LEFT (0xDA)
value VK_GAMEPAD_RIGHT_THUMBSTICK_RIGHT (0xD9)
value VK_GAMEPAD_RIGHT_THUMBSTICK_UP (0xD7)
value VK_GAMEPAD_RIGHT_TRIGGER (0xCA)
value VK_GAMEPAD_VIEW (0xD0)
value VK_GAMEPAD_X (0xC5)
value VK_GAMEPAD_Y (0xC6)
value VK_HANGEUL (0x15)
value VK_HANGUL (0x15)
value VK_HANJA (0x19)
value VK_HELP (0x2F)
value VK_HOME (0x24)
value VK_ICO_CLEAR (0xE6)
value VK_ICO_HELP (0xE3)
value VK_IME_OFF (0x1A)
value VK_IME_ON (0x16)
value VK_INSERT (0x2D)
value VK_JUNJA (0x17)
value VK_KANA (0x15)
value VK_KANJI (0x19)
value VK_LAUNCH_MAIL (0xB4)
value VK_LAUNCH_MEDIA_SELECT (0xB5)
value VK_LBUTTON (0x01)
value VK_LCONTROL (0xA2)
value VK_LEFT (0x25)
value VK_LMENU (0xA4)
value VK_LSHIFT (0xA0)
value VK_LWIN (0x5B)
value VK_MBUTTON (0x04)
value VK_MEDIA_NEXT_TRACK (0xB0)
value VK_MEDIA_PLAY_PAUSE (0xB3)
value VK_MEDIA_PREV_TRACK (0xB1)
value VK_MEDIA_STOP (0xB2)
value VK_MENU (0x12)
value VK_MODECHANGE (0x1F)
value VK_MULTIPLY (0x6A)
value VK_NAVIGATION_ACCEPT (0x8E)
value VK_NAVIGATION_CANCEL (0x8F)
value VK_NAVIGATION_DOWN (0x8B)
value VK_NAVIGATION_LEFT (0x8C)
value VK_NAVIGATION_MENU (0x89)
value VK_NAVIGATION_RIGHT (0x8D)
value VK_NAVIGATION_UP (0x8A)
value VK_NAVIGATION_VIEW (0x88)
value VK_NEXT (0x22)
value VK_NONAME (0xFC)
value VK_NONCONVERT (0x1D)
value VK_NUMLOCK (0x90)
value VK_OEM_ATTN (0xF0)
value VK_OEM_AUTO (0xF3)
value VK_OEM_AX (0xE1)
value VK_OEM_BACKTAB (0xF5)
value VK_OEM_CLEAR (0xFE)
value VK_OEM_COMMA (0xBC)
value VK_OEM_COPY (0xF2)
value VK_OEM_CUSEL (0xEF)
value VK_OEM_ENLW (0xF4)
value VK_OEM_FINISH (0xF1)
value VK_OEM_FJ_JISHO (0x92)
value VK_OEM_FJ_LOYA (0x95)
value VK_OEM_FJ_MASSHOU (0x93)
value VK_OEM_FJ_ROYA (0x96)
value VK_OEM_FJ_TOUROKU (0x94)
value VK_OEM_JUMP (0xEA)
value VK_OEM_MINUS (0xBD)
value VK_OEM_NEC_EQUAL (0x92)
value VK_OEM_PERIOD (0xBE)
value VK_OEM_PLUS (0xBB)
value VK_OEM_RESET (0xE9)
value VK_OEM_WSCTRL (0xEE)
value VK_PACKET (0xE7)
value VK_PAUSE (0x13)
value VK_PLAY (0xFA)
value VK_PRINT (0x2A)
value VK_PRIOR (0x21)
value VK_PROCESSKEY (0xE5)
value VK_RBUTTON (0x02)
value VK_RCONTROL (0xA3)
value VK_RETURN (0x0D)
value VK_RIGHT (0x27)
value VK_RMENU (0xA5)
value VK_RSHIFT (0xA1)
value VK_RWIN (0x5C)
value VK_SCROLL (0x91)
value VK_SELECT (0x29)
value VK_SEPARATOR (0x6C)
value VK_SHIFT (0x10)
value VK_SLEEP (0x5F)
value VK_SNAPSHOT (0x2C)
value VK_SPACE (0x20)
value VK_SUBTRACT (0x6D)
value VK_TAB (0x09)
value VK_UP (0x26)
value VK_VOLUME_DOWN (0xAE)
value VK_VOLUME_MUTE (0xAD)
value VK_VOLUME_UP (0xAF)
value VK_ZOOM (0xFB)
value VM_SAVED_STATE_DUMP_E_GUEST_MEMORY_NOT_FOUND (_HRESULT_TYPEDEF_(0xC0370501L))
value VM_SAVED_STATE_DUMP_E_INVALID_VP_STATE (_HRESULT_TYPEDEF_(0xC0370506L))
value VM_SAVED_STATE_DUMP_E_NESTED_VIRTUALIZATION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0xC0370503L))
value VM_SAVED_STATE_DUMP_E_NO_VP_FOUND_IN_PARTITION_STATE (_HRESULT_TYPEDEF_(0xC0370502L))
value VM_SAVED_STATE_DUMP_E_PARTITION_STATE_NOT_FOUND (_HRESULT_TYPEDEF_(0xC0370500L))
value VM_SAVED_STATE_DUMP_E_VA_NOT_MAPPED (_HRESULT_TYPEDEF_(0xC0370505L))
value VM_SAVED_STATE_DUMP_E_VP_VTL_NOT_ENABLED (_HRESULT_TYPEDEF_(0xC0370509L))
value VM_SAVED_STATE_DUMP_E_WINDOWS_KERNEL_IMAGE_NOT_FOUND (_HRESULT_TYPEDEF_(0xC0370504L))
value VOLUME_IS_DIRTY ((0x00000001))
value VOLUME_NAME_DOS (0x0)
value VOLUME_NAME_GUID (0x1)
value VOLUME_NAME_NONE (0x4)
value VOLUME_NAME_NT (0x2)
value VOLUME_SESSION_OPEN ((0x00000004))
value VOLUME_UPGRADE_SCHEDULED ((0x00000002))
value VOS_DOS (0x00010000L)
value VOS_NT (0x00040000L)
value VOS_UNKNOWN (0x00000000L)
value VOS_WINCE (0x00050000L)
value VOS__BASE (0x00000000L)
value VP_COMMAND_GET (0x0001)
value VP_COMMAND_SET (0x0002)
value VP_CP_CMD_ACTIVATE (0x0001)
value VP_CP_CMD_CHANGE (0x0004)
value VP_CP_CMD_DEACTIVATE (0x0002)
value VP_CP_TYPE_APS_TRIGGER (0x0001)
value VP_CP_TYPE_MACROVISION (0x0002)
value VP_FLAGS_BRIGHTNESS (0x0040)
value VP_FLAGS_CONTRAST (0x0080)
value VP_FLAGS_COPYPROTECT (0x0100)
value VP_FLAGS_FLICKER (0x0004)
value VP_FLAGS_MAX_UNSCALED (0x0010)
value VP_FLAGS_OVERSCAN (0x0008)
value VP_FLAGS_POSITION (0x0020)
value VP_FLAGS_TV_MODE (0x0001)
value VP_FLAGS_TV_STANDARD (0x0002)
value VP_MODE_TV_PLAYBACK (0x0002)
value VP_MODE_WIN_GRAPHICS (0x0001)
value VP_TV_STANDARD_NTSC_M (0x0001)
value VP_TV_STANDARD_NTSC_M_J (0x0002)
value VP_TV_STANDARD_PAL_B (0x0004)
value VP_TV_STANDARD_PAL_D (0x0008)
value VP_TV_STANDARD_PAL_G (0x00020000)
value VP_TV_STANDARD_PAL_H (0x0010)
value VP_TV_STANDARD_PAL_I (0x0020)
value VP_TV_STANDARD_PAL_M (0x0040)
value VP_TV_STANDARD_PAL_N (0x0080)
value VP_TV_STANDARD_SECAM_B (0x0100)
value VP_TV_STANDARD_SECAM_D (0x0200)
value VP_TV_STANDARD_SECAM_G (0x0400)
value VP_TV_STANDARD_SECAM_H (0x0800)
value VP_TV_STANDARD_SECAM_K (0x1000)
value VP_TV_STANDARD_SECAM_L (0x4000)
value VP_TV_STANDARD_WIN_VGA (0x8000)
value VREFRESH (116)
value VS_ALLOW_LATIN (0x0001)
value VS_FFI_FILEFLAGSMASK (0x0000003FL)
value VS_FFI_SIGNATURE (0xFEEF04BDL)
value VS_FFI_STRUCVERSION (0x00010000L)
value VS_FF_DEBUG (0x00000001L)
value VS_FF_INFOINFERRED (0x00000010L)
value VS_FF_PATCHED (0x00000004L)
value VS_FF_PRERELEASE (0x00000002L)
value VS_FF_PRIVATEBUILD (0x00000008L)
value VS_FF_SPECIALBUILD (0x00000020L)
value VS_FILE_INFO (RT_VERSION)
value VS_USER_DEFINED (100)
value VS_VERSION_INFO (1)
value VTA_BASELINE (TA_BASELINE)
value VTA_BOTTOM (TA_RIGHT)
value VTA_CENTER (TA_CENTER)
value VTA_LEFT (TA_BOTTOM)
value VTA_RIGHT (TA_TOP)
value VTA_TOP (TA_LEFT)
value VTDATEGRE_MAX (2958465)
value VTDATEGRE_MIN (-657434)
value VT_HARDTYPE (32768)
value WAIT_ABANDONED (((STATUS_ABANDONED_WAIT_0 ) + 0 ))
value WAIT_FAILED (((DWORD)0xFFFFFFFF))
value WAIT_IO_COMPLETION (STATUS_USER_APC)
value WAIT_TIMEOUT (258)
value WARNING_IPSEC_MM_POLICY_PRUNED (13024)
value WARNING_IPSEC_QM_POLICY_PRUNED (13025)
value WAVECAPS_LRVOLUME (0x0008)
value WAVECAPS_PITCH (0x0001)
value WAVECAPS_PLAYBACKRATE (0x0002)
value WAVECAPS_SAMPLEACCURATE (0x0020)
value WAVECAPS_SYNC (0x0010)
value WAVECAPS_VOLUME (0x0004)
value WAVERR_BADFORMAT ((WAVERR_BASE + 0))
value WAVERR_BASE (32)
value WAVERR_LASTERROR ((WAVERR_BASE + 3))
value WAVERR_STILLPLAYING ((WAVERR_BASE + 1))
value WAVERR_SYNC ((WAVERR_BASE + 3))
value WAVERR_UNPREPARED ((WAVERR_BASE + 2))
value WAVE_ALLOWSYNC (0x0002)
value WAVE_FORMAT_DIRECT (0x0008)
value WAVE_FORMAT_DIRECT_QUERY ((WAVE_FORMAT_QUERY | WAVE_FORMAT_DIRECT))
value WAVE_FORMAT_PCM (1)
value WAVE_FORMAT_QUERY (0x0001)
value WAVE_INVALIDFORMAT (0x00000000)
value WAVE_MAPPED (0x0004)
value WAVE_MAPPED_DEFAULT_COMMUNICATION_DEVICE (0x0010)
value WAVE_MAPPER (((UINT)-1))
value WA_ACTIVE (1)
value WA_CLICKACTIVE (2)
value WA_INACTIVE (0)
value WB_ISDELIMITER (2)
value WB_LEFT (0)
value WB_RIGHT (1)
value WC_COMPOSITECHECK (0x00000200)
value WC_DEFAULTCHAR (0x00000040)
value WC_DIALOG ((MAKEINTATOM(0x8002)))
value WC_DISCARDNS (0x00000010)
value WC_ERR_INVALID_CHARS (0x00000080)
value WC_NO_BEST_FIT_CHARS (0x00000400)
value WC_SEPCHARS (0x00000020)
value WDA_EXCLUDEFROMCAPTURE (0x00000011)
value WDA_MONITOR (0x00000001)
value WDA_NONE (0x00000000)
value WDK_NTDDI_VERSION (NTDDI_WIN10_NI)
value WDT_INPROC_CALL (( 0x48746457 ))
value WDT_REMOTE_CALL (( 0x52746457 ))
value WEB_E_INVALID_JSON_NUMBER (_HRESULT_TYPEDEF_(0x83750008L))
value WEB_E_INVALID_JSON_STRING (_HRESULT_TYPEDEF_(0x83750007L))
value WEB_E_INVALID_XML (_HRESULT_TYPEDEF_(0x83750002L))
value WEB_E_JSON_VALUE_NOT_FOUND (_HRESULT_TYPEDEF_(0x83750009L))
value WEB_E_MISSING_REQUIRED_ATTRIBUTE (_HRESULT_TYPEDEF_(0x83750004L))
value WEB_E_MISSING_REQUIRED_ELEMENT (_HRESULT_TYPEDEF_(0x83750003L))
value WEB_E_RESOURCE_TOO_LARGE (_HRESULT_TYPEDEF_(0x83750006L))
value WEB_E_UNEXPECTED_CONTENT (_HRESULT_TYPEDEF_(0x83750005L))
value WEB_E_UNSUPPORTED_FORMAT (_HRESULT_TYPEDEF_(0x83750001L))
value WEP_E_BUFFER_TOO_LARGE (_HRESULT_TYPEDEF_(0x88010009L))
value WEP_E_FIXED_DATA_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x88010002L))
value WEP_E_HARDWARE_NOT_COMPLIANT (_HRESULT_TYPEDEF_(0x88010003L))
value WEP_E_LOCK_NOT_CONFIGURED (_HRESULT_TYPEDEF_(0x88010004L))
value WEP_E_NOT_PROVISIONED_ON_ALL_VOLUMES (_HRESULT_TYPEDEF_(0x88010001L))
value WEP_E_NO_LICENSE (_HRESULT_TYPEDEF_(0x88010006L))
value WEP_E_OS_NOT_PROTECTED (_HRESULT_TYPEDEF_(0x88010007L))
value WEP_E_PROTECTION_SUSPENDED (_HRESULT_TYPEDEF_(0x88010005L))
value WEP_E_UNEXPECTED_FAIL (_HRESULT_TYPEDEF_(0x88010008L))
value WER_E_ALREADY_REPORTING (_HRESULT_TYPEDEF_(0x801B8004L))
value WER_E_CANCELED (_HRESULT_TYPEDEF_(0x801B8001L))
value WER_E_CRASH_FAILURE (_HRESULT_TYPEDEF_(0x801B8000L))
value WER_E_DUMP_THROTTLED (_HRESULT_TYPEDEF_(0x801B8005L))
value WER_E_INSUFFICIENT_CONSENT (_HRESULT_TYPEDEF_(0x801B8006L))
value WER_E_NETWORK_FAILURE (_HRESULT_TYPEDEF_(0x801B8002L))
value WER_E_NOT_INITIALIZED (_HRESULT_TYPEDEF_(0x801B8003L))
value WER_E_TOO_HEAVY (_HRESULT_TYPEDEF_(0x801B8007L))
value WER_S_ASSERT_CONTINUE (_HRESULT_TYPEDEF_(0x001B000AL))
value WER_S_DISABLED (_HRESULT_TYPEDEF_(0x001B0003L))
value WER_S_DISABLED_ARCHIVE (_HRESULT_TYPEDEF_(0x001B0006L))
value WER_S_DISABLED_QUEUE (_HRESULT_TYPEDEF_(0x001B0005L))
value WER_S_IGNORE_ALL_ASSERTS (_HRESULT_TYPEDEF_(0x001B0009L))
value WER_S_IGNORE_ASSERT_INSTANCE (_HRESULT_TYPEDEF_(0x001B0008L))
value WER_S_REPORT_ASYNC (_HRESULT_TYPEDEF_(0x001B0007L))
value WER_S_REPORT_DEBUG (_HRESULT_TYPEDEF_(0x001B0000L))
value WER_S_REPORT_QUEUED (_HRESULT_TYPEDEF_(0x001B0002L))
value WER_S_REPORT_UPLOADED (_HRESULT_TYPEDEF_(0x001B0001L))
value WER_S_REPORT_UPLOADED_CAB (_HRESULT_TYPEDEF_(0x001B000CL))
value WER_S_SUSPENDED_UPLOAD (_HRESULT_TYPEDEF_(0x001B0004L))
value WER_S_THROTTLED (_HRESULT_TYPEDEF_(0x001B000BL))
value WGL_FONT_LINES (0)
value WGL_FONT_POLYGONS (1)
value WGL_SWAPMULTIPLE_MAX (16)
value WGL_SWAP_MAIN_PLANE (0x00000001)
value WHDR_BEGINLOOP (0x00000004)
value WHDR_DONE (0x00000001)
value WHDR_ENDLOOP (0x00000008)
value WHDR_INQUEUE (0x00000010)
value WHDR_PREPARED (0x00000002)
value WHEEL_DELTA (120)
value WHEEL_PAGESCROLL ((UINT_MAX))
value WHITENESS ((DWORD)0x00FF0062)
value WHITEONBLACK (2)
value WHITE_BRUSH (0)
value WHITE_PEN (6)
value WHV_E_GPA_RANGE_NOT_FOUND (_HRESULT_TYPEDEF_(0x80370305L))
value WHV_E_INSUFFICIENT_BUFFER (_HRESULT_TYPEDEF_(0x80370301L))
value WHV_E_INVALID_PARTITION_CONFIG (_HRESULT_TYPEDEF_(0x80370304L))
value WHV_E_INVALID_VP_REGISTER_NAME (_HRESULT_TYPEDEF_(0x80370309L))
value WHV_E_INVALID_VP_STATE (_HRESULT_TYPEDEF_(0x80370308L))
value WHV_E_UNKNOWN_CAPABILITY (_HRESULT_TYPEDEF_(0x80370300L))
value WHV_E_UNKNOWN_PROPERTY (_HRESULT_TYPEDEF_(0x80370302L))
value WHV_E_UNSUPPORTED_HYPERVISOR_CONFIG (_HRESULT_TYPEDEF_(0x80370303L))
value WHV_E_UNSUPPORTED_PROCESSOR_CONFIG (_HRESULT_TYPEDEF_(0x80370310L))
value WHV_E_VP_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x80370306L))
value WHV_E_VP_DOES_NOT_EXIST (_HRESULT_TYPEDEF_(0x80370307L))
value WH_CALLWNDPROC (4)
value WH_CALLWNDPROCRET (12)
value WH_CBT (5)
value WH_DEBUG (9)
value WH_FOREGROUNDIDLE (11)
value WH_GETMESSAGE (3)
value WH_JOURNALPLAYBACK (1)
value WH_JOURNALRECORD (0)
value WH_KEYBOARD (2)
value WH_KEYBOARD_LL (13)
value WH_MAX (14)
value WH_MAXHOOK (WH_MAX)
value WH_MIN ((-1))
value WH_MINHOOK (WH_MIN)
value WH_MOUSE (7)
value WH_MOUSE_LL (14)
value WH_MSGFILTER ((-1))
value WH_SHELL (10)
value WH_SYSMSGFILTER (6)
value WIM_BOOT_NOT_OS_WIM ((0x00000000))
value WIM_BOOT_OS_WIM ((0x00000001))
value WIM_CLOSE (MM_WIM_CLOSE)
value WIM_DATA (MM_WIM_DATA)
value WIM_OPEN (MM_WIM_OPEN)
value WIM_PROVIDER_CURRENT_VERSION ((0x00000001))
value WIM_PROVIDER_EXTERNAL_FLAG_NOT_ACTIVE ((0x00000001))
value WIM_PROVIDER_EXTERNAL_FLAG_SUSPENDED ((0x00000002))
value WIM_PROVIDER_HASH_SIZE (20)
value WINABLEAPI (DECLSPEC_IMPORT)
value WINADVAPI (DECLSPEC_IMPORT)
value WINAPI_FAMILY (WINAPI_FAMILY_DESKTOP_APP)
value WINAPI_FAMILY_APP (WINAPI_FAMILY_PC_APP)
value WINAPI_FAMILY_DESKTOP_APP (100)
value WINAPI_FAMILY_GAMES (6)
value WINAPI_FAMILY_PC_APP (2)
value WINAPI_FAMILY_PHONE_APP (3)
value WINAPI_FAMILY_SERVER (5)
value WINAPI_FAMILY_SYSTEM (4)
value WINAPI_INLINE (WINAPI)
value WINAPI_PARTITION_PHONE (WINAPI_PARTITION_PHONE_APP)
value WINBASEAPI (DECLSPEC_IMPORT)
value WINCODEC_ERR_ALREADYLOCKED (_HRESULT_TYPEDEF_(0x88982F0DL))
value WINCODEC_ERR_BADHEADER (_HRESULT_TYPEDEF_(0x88982F61L))
value WINCODEC_ERR_BADIMAGE (_HRESULT_TYPEDEF_(0x88982F60L))
value WINCODEC_ERR_BADMETADATAHEADER (_HRESULT_TYPEDEF_(0x88982F63L))
value WINCODEC_ERR_BADSTREAMDATA (_HRESULT_TYPEDEF_(0x88982F70L))
value WINCODEC_ERR_CODECNOTHUMBNAIL (_HRESULT_TYPEDEF_(0x88982F44L))
value WINCODEC_ERR_CODECPRESENT (_HRESULT_TYPEDEF_(0x88982F43L))
value WINCODEC_ERR_CODECTOOMANYSCANLINES (_HRESULT_TYPEDEF_(0x88982F46L))
value WINCODEC_ERR_COMPONENTINITIALIZEFAILURE (_HRESULT_TYPEDEF_(0x88982F8BL))
value WINCODEC_ERR_COMPONENTNOTFOUND (_HRESULT_TYPEDEF_(0x88982F50L))
value WINCODEC_ERR_DUPLICATEMETADATAPRESENT (_HRESULT_TYPEDEF_(0x88982F8DL))
value WINCODEC_ERR_FRAMEMISSING (_HRESULT_TYPEDEF_(0x88982F62L))
value WINCODEC_ERR_IMAGESIZEOUTOFRANGE (_HRESULT_TYPEDEF_(0x88982F51L))
value WINCODEC_ERR_INSUFFICIENTBUFFER (_HRESULT_TYPEDEF_(0x88982F8CL))
value WINCODEC_ERR_INTERNALERROR (_HRESULT_TYPEDEF_(0x88982F48L))
value WINCODEC_ERR_INVALIDJPEGSCANINDEX (_HRESULT_TYPEDEF_(0x88982F96L))
value WINCODEC_ERR_INVALIDPROGRESSIVELEVEL (_HRESULT_TYPEDEF_(0x88982F95L))
value WINCODEC_ERR_INVALIDQUERYCHARACTER (_HRESULT_TYPEDEF_(0x88982F93L))
value WINCODEC_ERR_INVALIDQUERYREQUEST (_HRESULT_TYPEDEF_(0x88982F90L))
value WINCODEC_ERR_INVALIDREGISTRATION (_HRESULT_TYPEDEF_(0x88982F8AL))
value WINCODEC_ERR_NOTINITIALIZED (_HRESULT_TYPEDEF_(0x88982F0CL))
value WINCODEC_ERR_PALETTEUNAVAILABLE (_HRESULT_TYPEDEF_(0x88982F45L))
value WINCODEC_ERR_PROPERTYNOTFOUND (_HRESULT_TYPEDEF_(0x88982F40L))
value WINCODEC_ERR_PROPERTYNOTSUPPORTED (_HRESULT_TYPEDEF_(0x88982F41L))
value WINCODEC_ERR_PROPERTYSIZE (_HRESULT_TYPEDEF_(0x88982F42L))
value WINCODEC_ERR_PROPERTYUNEXPECTEDTYPE (_HRESULT_TYPEDEF_(0x88982F8EL))
value WINCODEC_ERR_REQUESTONLYVALIDATMETADATAROOT (_HRESULT_TYPEDEF_(0x88982F92L))
value WINCODEC_ERR_SOURCERECTDOESNOTMATCHDIMENSIONS (_HRESULT_TYPEDEF_(0x88982F49L))
value WINCODEC_ERR_STREAMNOTAVAILABLE (_HRESULT_TYPEDEF_(0x88982F73L))
value WINCODEC_ERR_STREAMREAD (_HRESULT_TYPEDEF_(0x88982F72L))
value WINCODEC_ERR_STREAMWRITE (_HRESULT_TYPEDEF_(0x88982F71L))
value WINCODEC_ERR_TOOMUCHMETADATA (_HRESULT_TYPEDEF_(0x88982F52L))
value WINCODEC_ERR_UNEXPECTEDMETADATATYPE (_HRESULT_TYPEDEF_(0x88982F91L))
value WINCODEC_ERR_UNEXPECTEDSIZE (_HRESULT_TYPEDEF_(0x88982F8FL))
value WINCODEC_ERR_UNKNOWNIMAGEFORMAT (_HRESULT_TYPEDEF_(0x88982F07L))
value WINCODEC_ERR_UNSUPPORTEDOPERATION (_HRESULT_TYPEDEF_(0x88982F81L))
value WINCODEC_ERR_UNSUPPORTEDPIXELFORMAT (_HRESULT_TYPEDEF_(0x88982F80L))
value WINCODEC_ERR_UNSUPPORTEDVERSION (_HRESULT_TYPEDEF_(0x88982F0BL))
value WINCODEC_ERR_VALUEOUTOFRANGE (_HRESULT_TYPEDEF_(0x88982F05L))
value WINCODEC_ERR_WRONGSTATE (_HRESULT_TYPEDEF_(0x88982F04L))
value WINCOMMCTRLAPI (DECLSPEC_IMPORT)
value WINCOMMDLGAPI (DECLSPEC_IMPORT)
value WINDEVQUERYAPI (DECLSPEC_IMPORT)
value WINDING (2)
value WINDOW_BUFFER_SIZE_EVENT (0x0004)
value WINEFS_SETUSERKEY_SET_CAPABILITIES (0x00000001)
value WINEVENT_INCONTEXT (0x0004)
value WINEVENT_OUTOFCONTEXT (0x0000)
value WINEVENT_SKIPOWNPROCESS (0x0002)
value WINEVENT_SKIPOWNTHREAD (0x0001)
value WINGDIAPI (DECLSPEC_IMPORT)
value WININETINFO_OPTION_LOCK_HANDLE (65534)
value WININET_E_ASYNC_THREAD_FAILED (_HRESULT_TYPEDEF_(0x80072F0FL))
value WININET_E_BAD_AUTO_PROXY_SCRIPT (_HRESULT_TYPEDEF_(0x80072F86L))
value WININET_E_BAD_OPTION_LENGTH (_HRESULT_TYPEDEF_(0x80072EEAL))
value WININET_E_BAD_REGISTRY_PARAMETER (_HRESULT_TYPEDEF_(0x80072EF6L))
value WININET_E_CANNOT_CONNECT (_HRESULT_TYPEDEF_(0x80072EFDL))
value WININET_E_CHG_POST_IS_NON_SECURE (_HRESULT_TYPEDEF_(0x80072F0AL))
value WININET_E_CLIENT_AUTH_CERT_NEEDED (_HRESULT_TYPEDEF_(0x80072F0CL))
value WININET_E_CLIENT_AUTH_NOT_SETUP (_HRESULT_TYPEDEF_(0x80072F0EL))
value WININET_E_CONNECTION_ABORTED (_HRESULT_TYPEDEF_(0x80072EFEL))
value WININET_E_CONNECTION_RESET (_HRESULT_TYPEDEF_(0x80072EFFL))
value WININET_E_COOKIE_DECLINED (_HRESULT_TYPEDEF_(0x80072F82L))
value WININET_E_COOKIE_NEEDS_CONFIRMATION (_HRESULT_TYPEDEF_(0x80072F81L))
value WININET_E_DECODING_FAILED (_HRESULT_TYPEDEF_(0x80072F8FL))
value WININET_E_DIALOG_PENDING (_HRESULT_TYPEDEF_(0x80072F11L))
value WININET_E_DISCONNECTED (_HRESULT_TYPEDEF_(0x80072F83L))
value WININET_E_DOWNLEVEL_SERVER (_HRESULT_TYPEDEF_(0x80072F77L))
value WININET_E_EXTENDED_ERROR (_HRESULT_TYPEDEF_(0x80072EE3L))
value WININET_E_FAILED_DUETOSECURITYCHECK (_HRESULT_TYPEDEF_(0x80072F8BL))
value WININET_E_FORCE_RETRY (_HRESULT_TYPEDEF_(0x80072F00L))
value WININET_E_HANDLE_EXISTS (_HRESULT_TYPEDEF_(0x80072F04L))
value WININET_E_HEADER_ALREADY_EXISTS (_HRESULT_TYPEDEF_(0x80072F7BL))
value WININET_E_HEADER_NOT_FOUND (_HRESULT_TYPEDEF_(0x80072F76L))
value WININET_E_HTTPS_HTTP_SUBMIT_REDIR (_HRESULT_TYPEDEF_(0x80072F14L))
value WININET_E_HTTPS_TO_HTTP_ON_REDIR (_HRESULT_TYPEDEF_(0x80072F08L))
value WININET_E_HTTP_TO_HTTPS_ON_REDIR (_HRESULT_TYPEDEF_(0x80072F07L))
value WININET_E_INCORRECT_FORMAT (_HRESULT_TYPEDEF_(0x80072EFBL))
value WININET_E_INCORRECT_HANDLE_STATE (_HRESULT_TYPEDEF_(0x80072EF3L))
value WININET_E_INCORRECT_HANDLE_TYPE (_HRESULT_TYPEDEF_(0x80072EF2L))
value WININET_E_INCORRECT_PASSWORD (_HRESULT_TYPEDEF_(0x80072EEEL))
value WININET_E_INCORRECT_USER_NAME (_HRESULT_TYPEDEF_(0x80072EEDL))
value WININET_E_INTERNAL_ERROR (_HRESULT_TYPEDEF_(0x80072EE4L))
value WININET_E_INVALID_CA (_HRESULT_TYPEDEF_(0x80072F0DL))
value WININET_E_INVALID_HEADER (_HRESULT_TYPEDEF_(0x80072F79L))
value WININET_E_INVALID_OPERATION (_HRESULT_TYPEDEF_(0x80072EF0L))
value WININET_E_INVALID_OPTION (_HRESULT_TYPEDEF_(0x80072EE9L))
value WININET_E_INVALID_PROXY_REQUEST (_HRESULT_TYPEDEF_(0x80072F01L))
value WININET_E_INVALID_QUERY_REQUEST (_HRESULT_TYPEDEF_(0x80072F7AL))
value WININET_E_INVALID_SERVER_RESPONSE (_HRESULT_TYPEDEF_(0x80072F78L))
value WININET_E_INVALID_URL (_HRESULT_TYPEDEF_(0x80072EE5L))
value WININET_E_ITEM_NOT_FOUND (_HRESULT_TYPEDEF_(0x80072EFCL))
value WININET_E_LOGIN_FAILURE (_HRESULT_TYPEDEF_(0x80072EEFL))
value WININET_E_LOGIN_FAILURE_DISPLAY_ENTITY_BODY (_HRESULT_TYPEDEF_(0x80072F8EL))
value WININET_E_MIXED_SECURITY (_HRESULT_TYPEDEF_(0x80072F09L))
value WININET_E_NAME_NOT_RESOLVED (_HRESULT_TYPEDEF_(0x80072EE7L))
value WININET_E_NEED_UI (_HRESULT_TYPEDEF_(0x80072F02L))
value WININET_E_NOT_INITIALIZED (_HRESULT_TYPEDEF_(0x80072F8CL))
value WININET_E_NOT_PROXY_REQUEST (_HRESULT_TYPEDEF_(0x80072EF4L))
value WININET_E_NOT_REDIRECTED (_HRESULT_TYPEDEF_(0x80072F80L))
value WININET_E_NO_CALLBACK (_HRESULT_TYPEDEF_(0x80072EF9L))
value WININET_E_NO_CONTEXT (_HRESULT_TYPEDEF_(0x80072EF8L))
value WININET_E_NO_DIRECT_ACCESS (_HRESULT_TYPEDEF_(0x80072EF7L))
value WININET_E_NO_NEW_CONTAINERS (_HRESULT_TYPEDEF_(0x80072F13L))
value WININET_E_OPERATION_CANCELLED (_HRESULT_TYPEDEF_(0x80072EF1L))
value WININET_E_OPTION_NOT_SETTABLE (_HRESULT_TYPEDEF_(0x80072EEBL))
value WININET_E_OUT_OF_HANDLES (_HRESULT_TYPEDEF_(0x80072EE1L))
value WININET_E_POST_IS_NON_SECURE (_HRESULT_TYPEDEF_(0x80072F0BL))
value WININET_E_PROTOCOL_NOT_FOUND (_HRESULT_TYPEDEF_(0x80072EE8L))
value WININET_E_PROXY_SERVER_UNREACHABLE (_HRESULT_TYPEDEF_(0x80072F85L))
value WININET_E_REDIRECT_FAILED (_HRESULT_TYPEDEF_(0x80072F7CL))
value WININET_E_REDIRECT_NEEDS_CONFIRMATION (_HRESULT_TYPEDEF_(0x80072F88L))
value WININET_E_REDIRECT_SCHEME_CHANGE (_HRESULT_TYPEDEF_(0x80072F10L))
value WININET_E_REGISTRY_VALUE_NOT_FOUND (_HRESULT_TYPEDEF_(0x80072EF5L))
value WININET_E_REQUEST_PENDING (_HRESULT_TYPEDEF_(0x80072EFAL))
value WININET_E_RETRY_DIALOG (_HRESULT_TYPEDEF_(0x80072F12L))
value WININET_E_SECURITY_CHANNEL_ERROR (_HRESULT_TYPEDEF_(0x80072F7DL))
value WININET_E_SEC_CERT_CN_INVALID (_HRESULT_TYPEDEF_(0x80072F06L))
value WININET_E_SEC_CERT_DATE_INVALID (_HRESULT_TYPEDEF_(0x80072F05L))
value WININET_E_SEC_CERT_ERRORS (_HRESULT_TYPEDEF_(0x80072F17L))
value WININET_E_SEC_CERT_REVOKED (_HRESULT_TYPEDEF_(0x80072F8AL))
value WININET_E_SEC_CERT_REV_FAILED (_HRESULT_TYPEDEF_(0x80072F19L))
value WININET_E_SEC_INVALID_CERT (_HRESULT_TYPEDEF_(0x80072F89L))
value WININET_E_SERVER_UNREACHABLE (_HRESULT_TYPEDEF_(0x80072F84L))
value WININET_E_SHUTDOWN (_HRESULT_TYPEDEF_(0x80072EECL))
value WININET_E_TCPIP_NOT_INSTALLED (_HRESULT_TYPEDEF_(0x80072F7FL))
value WININET_E_TIMEOUT (_HRESULT_TYPEDEF_(0x80072EE2L))
value WININET_E_UNABLE_TO_CACHE_FILE (_HRESULT_TYPEDEF_(0x80072F7EL))
value WININET_E_UNABLE_TO_DOWNLOAD_SCRIPT (_HRESULT_TYPEDEF_(0x80072F87L))
value WININET_E_UNRECOGNIZED_SCHEME (_HRESULT_TYPEDEF_(0x80072EE6L))
value WINML_ERR_INVALID_BINDING (_HRESULT_TYPEDEF_(0x88900002L))
value WINML_ERR_INVALID_DEVICE (_HRESULT_TYPEDEF_(0x88900001L))
value WINML_ERR_SIZE_MISMATCH (_HRESULT_TYPEDEF_(0x88900004L))
value WINML_ERR_VALUE_NOTFOUND (_HRESULT_TYPEDEF_(0x88900003L))
value WINMMAPI (DECLSPEC_IMPORT)
value WINNORMALIZEAPI (DECLSPEC_IMPORT)
value WINOLEAPI (EXTERN_C DECLSPEC_IMPORT HRESULT STDAPICALLTYPE)
value WINOLEAUTAPI (EXTERN_C DECLSPEC_IMPORT HRESULT STDAPICALLTYPE)
value WINPATHCCHAPI (WINBASEAPI)
value WINPERF_LOG_DEBUG (2)
value WINPERF_LOG_NONE (0)
value WINPERF_LOG_USER (1)
value WINPERF_LOG_VERBOSE (3)
value WINSHELLAPI (DECLSPEC_IMPORT)
value WINSOCK_API_LINKAGE (DECLSPEC_IMPORT)
value WINSPOOLAPI (DECLSPEC_IMPORT)
value WINSTA_ACCESSCLIPBOARD (0x0004L)
value WINSTA_ACCESSGLOBALATOMS (0x0020L)
value WINSTA_ALL_ACCESS ((WINSTA_ENUMDESKTOPS | WINSTA_READATTRIBUTES | WINSTA_ACCESSCLIPBOARD | WINSTA_CREATEDESKTOP | WINSTA_WRITEATTRIBUTES | WINSTA_ACCESSGLOBALATOMS | WINSTA_EXITWINDOWS | WINSTA_ENUMERATE | WINSTA_READSCREEN))
value WINSTA_CREATEDESKTOP (0x0008L)
value WINSTA_ENUMDESKTOPS (0x0001L)
value WINSTA_ENUMERATE (0x0100L)
value WINSTA_EXITWINDOWS (0x0040L)
value WINSTA_READATTRIBUTES (0x0002L)
value WINSTA_READSCREEN (0x0200L)
value WINSTA_WRITEATTRIBUTES (0x0010L)
value WINSTORAGEAPI (DECLSPEC_IMPORT)
value WINSWDEVICEAPI (DECLSPEC_IMPORT)
value WINUSERAPI (DECLSPEC_IMPORT)
value WINVER (_WIN32_WINNT)
value WIZ_BODYCX (184)
value WIZ_BODYX (92)
value WIZ_CXBMP (80)
value WIZ_CXDLG (276)
value WIZ_CYDLG (140)
value WMSZ_BOTTOM (6)
value WMSZ_BOTTOMLEFT (7)
value WMSZ_BOTTOMRIGHT (8)
value WMSZ_LEFT (1)
value WMSZ_RIGHT (2)
value WMSZ_TOP (3)
value WMSZ_TOPLEFT (4)
value WMSZ_TOPRIGHT (5)
value WM_ACTIVATE (0x0006)
value WM_ACTIVATEAPP (0x001C)
value WM_AFXFIRST (0x0360)
value WM_AFXLAST (0x037F)
value WM_APP (0x8000)
value WM_APPCOMMAND (0x0319)
value WM_ASKCBFORMATNAME (0x030C)
value WM_CANCELJOURNAL (0x004B)
value WM_CANCELMODE (0x001F)
value WM_CAPTURECHANGED (0x0215)
value WM_CHANGECBCHAIN (0x030D)
value WM_CHANGEUISTATE (0x0127)
value WM_CHAR (0x0102)
value WM_CHARTOITEM (0x002F)
value WM_CHILDACTIVATE (0x0022)
value WM_CHOOSEFONT_GETLOGFONT ((WM_USER + 1))
value WM_CHOOSEFONT_SETFLAGS ((WM_USER + 102))
value WM_CHOOSEFONT_SETLOGFONT ((WM_USER + 101))
value WM_CLEAR (0x0303)
value WM_CLIPBOARDUPDATE (0x031D)
value WM_CLOSE (0x0010)
value WM_COMMAND (0x0111)
value WM_COMMNOTIFY (0x0044)
value WM_COMPACTING (0x0041)
value WM_COMPAREITEM (0x0039)
value WM_CONTEXTMENU (0x007B)
value WM_COPY (0x0301)
value WM_COPYDATA (0x004A)
value WM_CREATE (0x0001)
value WM_CTLCOLORBTN (0x0135)
value WM_CTLCOLORDLG (0x0136)
value WM_CTLCOLOREDIT (0x0133)
value WM_CTLCOLORLISTBOX (0x0134)
value WM_CTLCOLORMSGBOX (0x0132)
value WM_CTLCOLORSCROLLBAR (0x0137)
value WM_CTLCOLORSTATIC (0x0138)
value WM_CUT (0x0300)
value WM_DDE_ACK ((WM_DDE_FIRST+4))
value WM_DDE_ADVISE ((WM_DDE_FIRST+2))
value WM_DDE_DATA ((WM_DDE_FIRST+5))
value WM_DDE_EXECUTE ((WM_DDE_FIRST+8))
value WM_DDE_FIRST (0x03E0)
value WM_DDE_INITIATE ((WM_DDE_FIRST))
value WM_DDE_LAST ((WM_DDE_FIRST+8))
value WM_DDE_POKE ((WM_DDE_FIRST+7))
value WM_DDE_REQUEST ((WM_DDE_FIRST+6))
value WM_DDE_TERMINATE ((WM_DDE_FIRST+1))
value WM_DDE_UNADVISE ((WM_DDE_FIRST+3))
value WM_DEADCHAR (0x0103)
value WM_DELETEITEM (0x002D)
value WM_DESTROY (0x0002)
value WM_DESTROYCLIPBOARD (0x0307)
value WM_DEVICECHANGE (0x0219)
value WM_DEVMODECHANGE (0x001B)
value WM_DISPLAYCHANGE (0x007E)
value WM_DPICHANGED (0x02E0)
value WM_DPICHANGED_AFTERPARENT (0x02E3)
value WM_DPICHANGED_BEFOREPARENT (0x02E2)
value WM_DRAWCLIPBOARD (0x0308)
value WM_DRAWITEM (0x002B)
value WM_DROPFILES (0x0233)
value WM_DWMCOLORIZATIONCOLORCHANGED (0x0320)
value WM_DWMCOMPOSITIONCHANGED (0x031E)
value WM_DWMNCRENDERINGCHANGED (0x031F)
value WM_DWMSENDICONICLIVEPREVIEWBITMAP (0x0326)
value WM_DWMSENDICONICTHUMBNAIL (0x0323)
value WM_DWMWINDOWMAXIMIZEDCHANGE (0x0321)
value WM_ENABLE (0x000A)
value WM_ENDSESSION (0x0016)
value WM_ENTERIDLE (0x0121)
value WM_ENTERMENULOOP (0x0211)
value WM_ENTERSIZEMOVE (0x0231)
value WM_ERASEBKGND (0x0014)
value WM_EXITMENULOOP (0x0212)
value WM_EXITSIZEMOVE (0x0232)
value WM_FONTCHANGE (0x001D)
value WM_GESTURE (0x0119)
value WM_GESTURENOTIFY (0x011A)
value WM_GETDLGCODE (0x0087)
value WM_GETDPISCALEDSIZE (0x02E4)
value WM_GETFONT (0x0031)
value WM_GETHOTKEY (0x0033)
value WM_GETICON (0x007F)
value WM_GETMINMAXINFO (0x0024)
value WM_GETOBJECT (0x003D)
value WM_GETTEXT (0x000D)
value WM_GETTEXTLENGTH (0x000E)
value WM_GETTITLEBARINFOEX (0x033F)
value WM_HANDHELDFIRST (0x0358)
value WM_HANDHELDLAST (0x035F)
value WM_HELP (0x0053)
value WM_HOTKEY (0x0312)
value WM_HSCROLL (0x0114)
value WM_HSCROLLCLIPBOARD (0x030E)
value WM_ICONERASEBKGND (0x0027)
value WM_IME_CHAR (0x0286)
value WM_IME_COMPOSITION (0x010F)
value WM_IME_COMPOSITIONFULL (0x0284)
value WM_IME_CONTROL (0x0283)
value WM_IME_ENDCOMPOSITION (0x010E)
value WM_IME_KEYDOWN (0x0290)
value WM_IME_KEYLAST (0x010F)
value WM_IME_KEYUP (0x0291)
value WM_IME_NOTIFY (0x0282)
value WM_IME_REQUEST (0x0288)
value WM_IME_SELECT (0x0285)
value WM_IME_SETCONTEXT (0x0281)
value WM_IME_STARTCOMPOSITION (0x010D)
value WM_INITDIALOG (0x0110)
value WM_INITMENU (0x0116)
value WM_INITMENUPOPUP (0x0117)
value WM_INPUT (0x00FF)
value WM_INPUTLANGCHANGE (0x0051)
value WM_INPUTLANGCHANGEREQUEST (0x0050)
value WM_INPUT_DEVICE_CHANGE (0x00FE)
value WM_KEYDOWN (0x0100)
value WM_KEYFIRST (0x0100)
value WM_KEYLAST (0x0109)
value WM_KEYUP (0x0101)
value WM_KILLFOCUS (0x0008)
value WM_LBUTTONDBLCLK (0x0203)
value WM_LBUTTONDOWN (0x0201)
value WM_LBUTTONUP (0x0202)
value WM_MBUTTONDBLCLK (0x0209)
value WM_MBUTTONDOWN (0x0207)
value WM_MBUTTONUP (0x0208)
value WM_MDIACTIVATE (0x0222)
value WM_MDICASCADE (0x0227)
value WM_MDICREATE (0x0220)
value WM_MDIDESTROY (0x0221)
value WM_MDIGETACTIVE (0x0229)
value WM_MDIICONARRANGE (0x0228)
value WM_MDIMAXIMIZE (0x0225)
value WM_MDINEXT (0x0224)
value WM_MDIREFRESHMENU (0x0234)
value WM_MDIRESTORE (0x0223)
value WM_MDISETMENU (0x0230)
value WM_MDITILE (0x0226)
value WM_MEASUREITEM (0x002C)
value WM_MENUCHAR (0x0120)
value WM_MENUCOMMAND (0x0126)
value WM_MENUDRAG (0x0123)
value WM_MENUGETOBJECT (0x0124)
value WM_MENURBUTTONUP (0x0122)
value WM_MENUSELECT (0x011F)
value WM_MOUSEACTIVATE (0x0021)
value WM_MOUSEFIRST (0x0200)
value WM_MOUSEHOVER (0x02A1)
value WM_MOUSEHWHEEL (0x020E)
value WM_MOUSELAST (0x020E)
value WM_MOUSELEAVE (0x02A3)
value WM_MOUSEMOVE (0x0200)
value WM_MOUSEWHEEL (0x020A)
value WM_MOVE (0x0003)
value WM_MOVING (0x0216)
value WM_NCACTIVATE (0x0086)
value WM_NCCALCSIZE (0x0083)
value WM_NCCREATE (0x0081)
value WM_NCDESTROY (0x0082)
value WM_NCHITTEST (0x0084)
value WM_NCLBUTTONDBLCLK (0x00A3)
value WM_NCLBUTTONDOWN (0x00A1)
value WM_NCLBUTTONUP (0x00A2)
value WM_NCMBUTTONDBLCLK (0x00A9)
value WM_NCMBUTTONDOWN (0x00A7)
value WM_NCMBUTTONUP (0x00A8)
value WM_NCMOUSEHOVER (0x02A0)
value WM_NCMOUSELEAVE (0x02A2)
value WM_NCMOUSEMOVE (0x00A0)
value WM_NCPAINT (0x0085)
value WM_NCPOINTERDOWN (0x0242)
value WM_NCPOINTERUP (0x0243)
value WM_NCPOINTERUPDATE (0x0241)
value WM_NCRBUTTONDBLCLK (0x00A6)
value WM_NCRBUTTONDOWN (0x00A4)
value WM_NCRBUTTONUP (0x00A5)
value WM_NCXBUTTONDBLCLK (0x00AD)
value WM_NCXBUTTONDOWN (0x00AB)
value WM_NCXBUTTONUP (0x00AC)
value WM_NEXTDLGCTL (0x0028)
value WM_NEXTMENU (0x0213)
value WM_NOTIFY (0x004E)
value WM_NOTIFYFORMAT (0x0055)
value WM_NULL (0x0000)
value WM_PAINT (0x000F)
value WM_PAINTCLIPBOARD (0x0309)
value WM_PAINTICON (0x0026)
value WM_PALETTECHANGED (0x0311)
value WM_PALETTEISCHANGING (0x0310)
value WM_PARENTNOTIFY (0x0210)
value WM_PASTE (0x0302)
value WM_PENWINFIRST (0x0380)
value WM_PENWINLAST (0x038F)
value WM_POINTERACTIVATE (0x024B)
value WM_POINTERCAPTURECHANGED (0x024C)
value WM_POINTERDEVICECHANGE (0x238)
value WM_POINTERDEVICEINRANGE (0x239)
value WM_POINTERDEVICEOUTOFRANGE (0x23A)
value WM_POINTERDOWN (0x0246)
value WM_POINTERENTER (0x0249)
value WM_POINTERHWHEEL (0x024F)
value WM_POINTERLEAVE (0x024A)
value WM_POINTERROUTEDAWAY (0x0252)
value WM_POINTERROUTEDRELEASED (0x0253)
value WM_POINTERROUTEDTO (0x0251)
value WM_POINTERUP (0x0247)
value WM_POINTERUPDATE (0x0245)
value WM_POINTERWHEEL (0x024E)
value WM_POWER (0x0048)
value WM_POWERBROADCAST (0x0218)
value WM_PRINT (0x0317)
value WM_PRINTCLIENT (0x0318)
value WM_PSD_ENVSTAMPRECT ((WM_USER+5))
value WM_PSD_FULLPAGERECT ((WM_USER+1))
value WM_PSD_GREEKTEXTRECT ((WM_USER+4))
value WM_PSD_MARGINRECT ((WM_USER+3))
value WM_PSD_MINMARGINRECT ((WM_USER+2))
value WM_PSD_PAGESETUPDLG ((WM_USER ))
value WM_PSD_YAFULLPAGERECT ((WM_USER+6))
value WM_QUERYDRAGICON (0x0037)
value WM_QUERYENDSESSION (0x0011)
value WM_QUERYNEWPALETTE (0x030F)
value WM_QUERYOPEN (0x0013)
value WM_QUERYUISTATE (0x0129)
value WM_QUEUESYNC (0x0023)
value WM_QUIT (0x0012)
value WM_RBUTTONDBLCLK (0x0206)
value WM_RBUTTONDOWN (0x0204)
value WM_RBUTTONUP (0x0205)
value WM_RENDERALLFORMATS (0x0306)
value WM_RENDERFORMAT (0x0305)
value WM_SETCURSOR (0x0020)
value WM_SETFOCUS (0x0007)
value WM_SETFONT (0x0030)
value WM_SETHOTKEY (0x0032)
value WM_SETICON (0x0080)
value WM_SETREDRAW (0x000B)
value WM_SETTEXT (0x000C)
value WM_SETTINGCHANGE (WM_WININICHANGE)
value WM_SHOWWINDOW (0x0018)
value WM_SIZE (0x0005)
value WM_SIZECLIPBOARD (0x030B)
value WM_SIZING (0x0214)
value WM_SPOOLERSTATUS (0x002A)
value WM_STYLECHANGED (0x007D)
value WM_STYLECHANGING (0x007C)
value WM_SYNCPAINT (0x0088)
value WM_SYSCHAR (0x0106)
value WM_SYSCOLORCHANGE (0x0015)
value WM_SYSCOMMAND (0x0112)
value WM_SYSDEADCHAR (0x0107)
value WM_SYSKEYDOWN (0x0104)
value WM_SYSKEYUP (0x0105)
value WM_TABLET_FIRST (0x02c0)
value WM_TABLET_LAST (0x02df)
value WM_TCARD (0x0052)
value WM_THEMECHANGED (0x031A)
value WM_TIMECHANGE (0x001E)
value WM_TIMER (0x0113)
value WM_TOOLTIPDISMISS (0x0345)
value WM_TOUCH (0x0240)
value WM_TOUCHHITTESTING (0x024D)
value WM_UNDO (0x0304)
value WM_UNICHAR (0x0109)
value WM_UNINITMENUPOPUP (0x0125)
value WM_UPDATEUISTATE (0x0128)
value WM_USER (0x0400)
value WM_USERCHANGED (0x0054)
value WM_VKEYTOITEM (0x002E)
value WM_VSCROLL (0x0115)
value WM_VSCROLLCLIPBOARD (0x030A)
value WM_WINDOWPOSCHANGED (0x0047)
value WM_WINDOWPOSCHANGING (0x0046)
value WM_WININICHANGE (0x001A)
value WM_WTSSESSION_CHANGE (0x02B1)
value WM_XBUTTONDBLCLK (0x020D)
value WM_XBUTTONDOWN (0x020B)
value WM_XBUTTONUP (0x020C)
value WNCON_DYNAMIC (0x00000008)
value WNCON_FORNETCARD (0x00000001)
value WNCON_NOTROUTED (0x00000002)
value WNCON_SLOWLINK (0x00000004)
value WNFMT_ABBREVIATED (0x02)
value WNFMT_CONNECTION (0x20)
value WNFMT_INENUM (0x10)
value WNFMT_MULTILINE (0x01)
value WNNC_CRED_MANAGER (0xFFFF0000)
value WNNC_NET_APPLETALK (0x00130000)
value WNNC_NET_AURISTOR_FS (0x00460000)
value WNNC_NET_AVID (0x001A0000)
value WNNC_NET_BMC (0x00180000)
value WNNC_NET_BWNFS (0x00100000)
value WNNC_NET_CLEARCASE (0x00160000)
value WNNC_NET_COGENT (0x00110000)
value WNNC_NET_CSC (0x00260000)
value WNNC_NET_DAV (0x002E0000)
value WNNC_NET_DCE (0x00190000)
value WNNC_NET_DECORB (0x00200000)
value WNNC_NET_DFS (0x003B0000)
value WNNC_NET_DISTINCT (0x00230000)
value WNNC_NET_DOCUSHARE (0x00450000)
value WNNC_NET_DOCUSPACE (0x001B0000)
value WNNC_NET_DRIVEONWEB (0x003E0000)
value WNNC_NET_EXIFS (0x002D0000)
value WNNC_NET_EXTENDNET (0x00290000)
value WNNC_NET_FARALLON (0x00120000)
value WNNC_NET_FJ_REDIR (0x00220000)
value WNNC_NET_FOXBAT (0x002B0000)
value WNNC_NET_FRONTIER (0x00170000)
value WNNC_NET_FTP_NFS (0x000C0000)
value WNNC_NET_GOOGLE (0x00430000)
value WNNC_NET_HOB_NFS (0x00320000)
value WNNC_NET_IBMAL (0x00340000)
value WNNC_NET_INTERGRAPH (0x00140000)
value WNNC_NET_KNOWARE (0x002F0000)
value WNNC_NET_KWNP (0x003C0000)
value WNNC_NET_LANMAN (WNNC_NET_SMB)
value WNNC_NET_LANSTEP (0x00080000)
value WNNC_NET_LANTASTIC (0x000A0000)
value WNNC_NET_LIFENET (0x000E0000)
value WNNC_NET_LOCK (0x00350000)
value WNNC_NET_LOCUS (0x00060000)
value WNNC_NET_MANGOSOFT (0x001C0000)
value WNNC_NET_MASFAX (0x00310000)
value WNNC_NET_MFILES (0x00410000)
value WNNC_NET_MSNET (0x00010000)
value WNNC_NET_MS_NFS (0x00420000)
value WNNC_NET_NDFS (0x00440000)
value WNNC_NET_NETWARE (0x00030000)
value WNNC_NET_OBJECT_DIRE (0x00300000)
value WNNC_NET_OPENAFS (0x00390000)
value WNNC_NET_PATHWORKS (0x000D0000)
value WNNC_NET_POWERLAN (0x000F0000)
value WNNC_NET_PROTSTOR (0x00210000)
value WNNC_NET_QUINCY (0x00380000)
value WNNC_NET_RSFX (0x00400000)
value WNNC_NET_SECUREAGENT (0x00470000)
value WNNC_NET_SERNET (0x001D0000)
value WNNC_NET_SHIVA (0x00330000)
value WNNC_NET_SMB (0x00020000)
value WNNC_NET_SRT (0x00370000)
value WNNC_NET_STAC (0x002A0000)
value WNNC_NET_SUN_PC_NFS (0x00070000)
value WNNC_NET_SYMFONET (0x00150000)
value WNNC_NET_TERMSRV (0x00360000)
value WNNC_NET_TWINS (0x00240000)
value WNNC_NET_VINES (0x00040000)
value WNNC_NET_VMWARE (0x003F0000)
value WNNC_NET_YAHOO (0x002C0000)
value WNNC_NET_ZENWORKS (0x003D0000)
value WN_ACCESS_DENIED (ERROR_ACCESS_DENIED)
value WN_ALREADY_CONNECTED (ERROR_ALREADY_ASSIGNED)
value WN_BAD_DEV_TYPE (ERROR_BAD_DEV_TYPE)
value WN_BAD_HANDLE (ERROR_INVALID_HANDLE)
value WN_BAD_LEVEL (ERROR_INVALID_LEVEL)
value WN_BAD_LOCALNAME (ERROR_BAD_DEVICE)
value WN_BAD_NETNAME (ERROR_BAD_NET_NAME)
value WN_BAD_PASSWORD (ERROR_INVALID_PASSWORD)
value WN_BAD_POINTER (ERROR_INVALID_ADDRESS)
value WN_BAD_PROFILE (ERROR_BAD_PROFILE)
value WN_BAD_PROVIDER (ERROR_BAD_PROVIDER)
value WN_BAD_USER (ERROR_BAD_USERNAME)
value WN_BAD_VALUE (ERROR_INVALID_PARAMETER)
value WN_CANCEL (ERROR_CANCELLED)
value WN_CANNOT_OPEN_PROFILE (ERROR_CANNOT_OPEN_PROFILE)
value WN_CONNECTED_OTHER_PASSWORD (ERROR_CONNECTED_OTHER_PASSWORD)
value WN_CONNECTED_OTHER_PASSWORD_DEFAULT (ERROR_CONNECTED_OTHER_PASSWORD_DEFAULT)
value WN_CONNECTION_CLOSED (ERROR_CONNECTION_UNAVAIL)
value WN_DEVICE_ALREADY_REMEMBERED (ERROR_DEVICE_ALREADY_REMEMBERED)
value WN_DEVICE_ERROR (ERROR_GEN_FAILURE)
value WN_DEVICE_IN_USE (ERROR_DEVICE_IN_USE)
value WN_EXTENDED_ERROR (ERROR_EXTENDED_ERROR)
value WN_FUNCTION_BUSY (ERROR_BUSY)
value WN_MORE_DATA (ERROR_MORE_DATA)
value WN_NET_ERROR (ERROR_UNEXP_NET_ERR)
value WN_NOT_AUTHENTICATED (ERROR_NOT_AUTHENTICATED)
value WN_NOT_CONNECTED (ERROR_NOT_CONNECTED)
value WN_NOT_CONTAINER (ERROR_NOT_CONTAINER)
value WN_NOT_INITIALIZING (ERROR_ALREADY_INITIALIZED)
value WN_NOT_LOGGED_ON (ERROR_NOT_LOGGED_ON)
value WN_NOT_SUPPORTED (ERROR_NOT_SUPPORTED)
value WN_NOT_VALIDATED (ERROR_NO_LOGON_SERVERS)
value WN_NO_ERROR (NO_ERROR)
value WN_NO_MORE_DEVICES (ERROR_NO_MORE_DEVICES)
value WN_NO_MORE_ENTRIES (ERROR_NO_MORE_ITEMS)
value WN_NO_NETWORK (ERROR_NO_NETWORK)
value WN_NO_NET_OR_BAD_PATH (ERROR_NO_NET_OR_BAD_PATH)
value WN_OPEN_FILES (ERROR_OPEN_FILES)
value WN_OUT_OF_MEMORY (ERROR_NOT_ENOUGH_MEMORY)
value WN_RETRY (ERROR_RETRY)
value WN_SUCCESS (NO_ERROR)
value WN_WINDOWS_ERROR (ERROR_UNEXP_NET_ERR)
value WOF_CURRENT_VERSION ((0x00000001))
value WOF_PROVIDER_CLOUD ((0x00000003))
value WOF_PROVIDER_FILE ((0x00000002))
value WOF_PROVIDER_WIM ((0x00000001))
value WOM_CLOSE (MM_WOM_CLOSE)
value WOM_DONE (MM_WOM_DONE)
value WOM_OPEN (MM_WOM_OPEN)
value WPF_ASYNCWINDOWPLACEMENT (0x0004)
value WPF_RESTORETOMAXIMIZED (0x0002)
value WPF_SETMINPOSITION (0x0001)
value WPN_E_ACCESS_DENIED (_HRESULT_TYPEDEF_(0x803E0117L))
value WPN_E_ALL_URL_NOT_COMPLETED (_HRESULT_TYPEDEF_(0x803E0203L))
value WPN_E_CALLBACK_ALREADY_REGISTERED (_HRESULT_TYPEDEF_(0x803E0206L))
value WPN_E_CHANNEL_CLOSED (_HRESULT_TYPEDEF_(0x803E0100L))
value WPN_E_CHANNEL_REQUEST_NOT_COMPLETE (_HRESULT_TYPEDEF_(0x803E0101L))
value WPN_E_CLOUD_AUTH_UNAVAILABLE (_HRESULT_TYPEDEF_(0x803E011AL))
value WPN_E_CLOUD_DISABLED (_HRESULT_TYPEDEF_(0x803E0109L))
value WPN_E_CLOUD_DISABLED_FOR_APP (_HRESULT_TYPEDEF_(0x803E020BL))
value WPN_E_CLOUD_INCAPABLE (_HRESULT_TYPEDEF_(0x803E0110L))
value WPN_E_CLOUD_SERVICE_UNAVAILABLE (_HRESULT_TYPEDEF_(0x803E011BL))
value WPN_E_DEV_ID_SIZE (_HRESULT_TYPEDEF_(0x803E0120L))
value WPN_E_DUPLICATE_CHANNEL (_HRESULT_TYPEDEF_(0x803E0104L))
value WPN_E_DUPLICATE_REGISTRATION (_HRESULT_TYPEDEF_(0x803E0118L))
value WPN_E_FAILED_LOCK_SCREEN_UPDATE_INTIALIZATION (_HRESULT_TYPEDEF_(0x803E011CL))
value WPN_E_GROUP_ALPHANUMERIC (_HRESULT_TYPEDEF_(0x803E020AL))
value WPN_E_GROUP_SIZE (_HRESULT_TYPEDEF_(0x803E0209L))
value WPN_E_IMAGE_NOT_FOUND_IN_CACHE (_HRESULT_TYPEDEF_(0x803E0202L))
value WPN_E_INTERNET_INCAPABLE (_HRESULT_TYPEDEF_(0x803E0113L))
value WPN_E_INVALID_APP (_HRESULT_TYPEDEF_(0x803E0102L))
value WPN_E_INVALID_CLOUD_IMAGE (_HRESULT_TYPEDEF_(0x803E0204L))
value WPN_E_INVALID_HTTP_STATUS_CODE (_HRESULT_TYPEDEF_(0x803E012BL))
value WPN_E_NOTIFICATION_DISABLED (_HRESULT_TYPEDEF_(0x803E0111L))
value WPN_E_NOTIFICATION_HIDDEN (_HRESULT_TYPEDEF_(0x803E0107L))
value WPN_E_NOTIFICATION_ID_MATCHED (_HRESULT_TYPEDEF_(0x803E0205L))
value WPN_E_NOTIFICATION_INCAPABLE (_HRESULT_TYPEDEF_(0x803E0112L))
value WPN_E_NOTIFICATION_NOT_POSTED (_HRESULT_TYPEDEF_(0x803E0108L))
value WPN_E_NOTIFICATION_POSTED (_HRESULT_TYPEDEF_(0x803E0106L))
value WPN_E_NOTIFICATION_SIZE (_HRESULT_TYPEDEF_(0x803E0115L))
value WPN_E_NOTIFICATION_TYPE_DISABLED (_HRESULT_TYPEDEF_(0x803E0114L))
value WPN_E_OUTSTANDING_CHANNEL_REQUEST (_HRESULT_TYPEDEF_(0x803E0103L))
value WPN_E_OUT_OF_SESSION (_HRESULT_TYPEDEF_(0x803E0200L))
value WPN_E_PLATFORM_UNAVAILABLE (_HRESULT_TYPEDEF_(0x803E0105L))
value WPN_E_POWER_SAVE (_HRESULT_TYPEDEF_(0x803E0201L))
value WPN_E_PUSH_NOTIFICATION_INCAPABLE (_HRESULT_TYPEDEF_(0x803E0119L))
value WPN_E_STORAGE_LOCKED (_HRESULT_TYPEDEF_(0x803E0208L))
value WPN_E_TAG_ALPHANUMERIC (_HRESULT_TYPEDEF_(0x803E012AL))
value WPN_E_TAG_SIZE (_HRESULT_TYPEDEF_(0x803E0116L))
value WPN_E_TOAST_NOTIFICATION_DROPPED (_HRESULT_TYPEDEF_(0x803E0207L))
value WRITE_COMPRESSION_INFO_VALID (0x00000010)
value WRITE_DAC ((0x00040000L))
value WRITE_NV_MEMORY_FLAG_FLUSH ((0x00000001))
value WRITE_NV_MEMORY_FLAG_NON_TEMPORAL ((0x00000002))
value WRITE_NV_MEMORY_FLAG_NO_DRAIN ((0x00000100))
value WRITE_NV_MEMORY_FLAG_PERSIST ((WRITE_NV_MEMORY_FLAG_FLUSH | WRITE_NV_MEMORY_FLAG_NON_TEMPORAL))
value WRITE_OWNER ((0x00080000L))
value WRITE_RESTRICTED (0x8)
value WRITE_WATCH_FLAG_RESET (0x01)
value WSAAPI (FAR PASCAL)
value WSABASEERR (10000)
value WSADESCRIPTION_LEN (256)
value WSAEACCES (10013)
value WSAEADDRINUSE (10048)
value WSAEADDRNOTAVAIL (10049)
value WSAEAFNOSUPPORT (10047)
value WSAEALREADY (10037)
value WSAEBADF (10009)
value WSAECANCELLED (10103)
value WSAECONNABORTED (10053)
value WSAECONNREFUSED (10061)
value WSAECONNRESET (10054)
value WSAEDESTADDRREQ (10039)
value WSAEDISCON (10101)
value WSAEDQUOT (10069)
value WSAEFAULT (10014)
value WSAEHOSTDOWN (10064)
value WSAEHOSTUNREACH (10065)
value WSAEINPROGRESS (10036)
value WSAEINTR (10004)
value WSAEINVAL (10022)
value WSAEINVALIDPROCTABLE (10104)
value WSAEINVALIDPROVIDER (10105)
value WSAEISCONN (10056)
value WSAELOOP (10062)
value WSAEMFILE (10024)
value WSAEMSGSIZE (10040)
value WSAENAMETOOLONG (10063)
value WSAENETDOWN (10050)
value WSAENETRESET (10052)
value WSAENETUNREACH (10051)
value WSAENOBUFS (10055)
value WSAENOMORE (10102)
value WSAENOPROTOOPT (10042)
value WSAENOTCONN (10057)
value WSAENOTEMPTY (10066)
value WSAENOTSOCK (10038)
value WSAEOPNOTSUPP (10045)
value WSAEPFNOSUPPORT (10046)
value WSAEPROCLIM (10067)
value WSAEPROTONOSUPPORT (10043)
value WSAEPROTOTYPE (10041)
value WSAEPROVIDERFAILEDINIT (10106)
value WSAEREFUSED (10112)
value WSAEREMOTE (10071)
value WSAESHUTDOWN (10058)
value WSAESOCKTNOSUPPORT (10044)
value WSAESTALE (10070)
value WSAETIMEDOUT (10060)
value WSAETOOMANYREFS (10059)
value WSAEUSERS (10068)
value WSAEVENT (HANDLE)
value WSAEWOULDBLOCK (10035)
value WSAHOST_NOT_FOUND (11001)
value WSANOTINITIALISED (10093)
value WSANO_ADDRESS (WSANO_DATA)
value WSANO_DATA (11004)
value WSANO_RECOVERY (11003)
value WSAOVERLAPPED (OVERLAPPED)
value WSAPROTOCOL_LEN (255)
value WSASERVICE_NOT_FOUND (10108)
value WSASYSCALLFAILURE (10107)
value WSASYSNOTREADY (10091)
value WSASYS_STATUS_LEN (128)
value WSATRY_AGAIN (11002)
value WSATYPE_NOT_FOUND (10109)
value WSAVERNOTSUPPORTED (10092)
value WSA_E_CANCELLED (10111)
value WSA_E_NO_MORE (10110)
value WSA_FLAG_ACCESS_SYSTEM_SECURITY (0x40)
value WSA_FLAG_MULTIPOINT_C_LEAF (0x04)
value WSA_FLAG_MULTIPOINT_C_ROOT (0x02)
value WSA_FLAG_MULTIPOINT_D_LEAF (0x10)
value WSA_FLAG_MULTIPOINT_D_ROOT (0x08)
value WSA_FLAG_NO_HANDLE_INHERIT (0x80)
value WSA_FLAG_OVERLAPPED (0x01)
value WSA_FLAG_REGISTERED_IO (0x100)
value WSA_INFINITE ((INFINITE))
value WSA_INVALID_EVENT (((WSAEVENT)NULL))
value WSA_INVALID_HANDLE ((ERROR_INVALID_HANDLE))
value WSA_INVALID_PARAMETER ((ERROR_INVALID_PARAMETER))
value WSA_IO_INCOMPLETE ((ERROR_IO_INCOMPLETE))
value WSA_IO_PENDING ((ERROR_IO_PENDING))
value WSA_IPSEC_NAME_POLICY_ERROR (11033)
value WSA_MAXIMUM_WAIT_EVENTS ((MAXIMUM_WAIT_OBJECTS))
value WSA_NOT_ENOUGH_MEMORY ((ERROR_NOT_ENOUGH_MEMORY))
value WSA_OPERATION_ABORTED ((ERROR_OPERATION_ABORTED))
value WSA_QOS_ADMISSION_FAILURE (11010)
value WSA_QOS_BAD_OBJECT (11013)
value WSA_QOS_BAD_STYLE (11012)
value WSA_QOS_EFILTERCOUNT (11021)
value WSA_QOS_EFILTERSTYLE (11019)
value WSA_QOS_EFILTERTYPE (11020)
value WSA_QOS_EFLOWCOUNT (11023)
value WSA_QOS_EFLOWDESC (11026)
value WSA_QOS_EFLOWSPEC (11017)
value WSA_QOS_EOBJLENGTH (11022)
value WSA_QOS_EPOLICYOBJ (11025)
value WSA_QOS_EPROVSPECBUF (11018)
value WSA_QOS_EPSFILTERSPEC (11028)
value WSA_QOS_EPSFLOWSPEC (11027)
value WSA_QOS_ESDMODEOBJ (11029)
value WSA_QOS_ESERVICETYPE (11016)
value WSA_QOS_ESHAPERATEOBJ (11030)
value WSA_QOS_EUNKOWNPSOBJ (11024)
value WSA_QOS_GENERIC_ERROR (11015)
value WSA_QOS_NO_RECEIVERS (11008)
value WSA_QOS_NO_SENDERS (11007)
value WSA_QOS_POLICY_FAILURE (11011)
value WSA_QOS_RECEIVERS (11005)
value WSA_QOS_REQUEST_CONFIRMED (11009)
value WSA_QOS_RESERVED_PETYPE (11031)
value WSA_QOS_SENDERS (11006)
value WSA_QOS_TRAFFIC_CTRL_ERROR (11014)
value WSA_SECURE_HOST_NOT_FOUND (11032)
value WSA_WAIT_FAILED ((WAIT_FAILED))
value WSA_WAIT_IO_COMPLETION ((WAIT_IO_COMPLETION))
value WSA_WAIT_TIMEOUT ((WAIT_TIMEOUT))
value WSF_VISIBLE (0x0001L)
value WSK_SO_BASE (0x4000)
value WS_ACTIVECAPTION (0x0001)
value WS_BORDER (0x00800000L)
value WS_CAPTION (0x00C00000L)
value WS_CHILD (0x40000000L)
value WS_CHILDWINDOW ((WS_CHILD))
value WS_CLIPCHILDREN (0x02000000L)
value WS_CLIPSIBLINGS (0x04000000L)
value WS_DISABLED (0x08000000L)
value WS_DLGFRAME (0x00400000L)
value WS_EX_ACCEPTFILES (0x00000010L)
value WS_EX_APPWINDOW (0x00040000L)
value WS_EX_CLIENTEDGE (0x00000200L)
value WS_EX_COMPOSITED (0x02000000L)
value WS_EX_CONTEXTHELP (0x00000400L)
value WS_EX_CONTROLPARENT (0x00010000L)
value WS_EX_DLGMODALFRAME (0x00000001L)
value WS_EX_LAYERED (0x00080000)
value WS_EX_LAYOUTRTL (0x00400000L)
value WS_EX_LEFT (0x00000000L)
value WS_EX_LEFTSCROLLBAR (0x00004000L)
value WS_EX_LTRREADING (0x00000000L)
value WS_EX_MDICHILD (0x00000040L)
value WS_EX_NOACTIVATE (0x08000000L)
value WS_EX_NOINHERITLAYOUT (0x00100000L)
value WS_EX_NOPARENTNOTIFY (0x00000004L)
value WS_EX_NOREDIRECTIONBITMAP (0x00200000L)
value WS_EX_OVERLAPPEDWINDOW ((WS_EX_WINDOWEDGE | WS_EX_CLIENTEDGE))
value WS_EX_PALETTEWINDOW ((WS_EX_WINDOWEDGE | WS_EX_TOOLWINDOW | WS_EX_TOPMOST))
value WS_EX_RIGHT (0x00001000L)
value WS_EX_RIGHTSCROLLBAR (0x00000000L)
value WS_EX_RTLREADING (0x00002000L)
value WS_EX_STATICEDGE (0x00020000L)
value WS_EX_TOOLWINDOW (0x00000080L)
value WS_EX_TOPMOST (0x00000008L)
value WS_EX_TRANSPARENT (0x00000020L)
value WS_EX_WINDOWEDGE (0x00000100L)
value WS_E_ADDRESS_IN_USE (_HRESULT_TYPEDEF_(0x803D000BL))
value WS_E_ADDRESS_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x803D000CL))
value WS_E_ENDPOINT_ACCESS_DENIED (_HRESULT_TYPEDEF_(0x803D0005L))
value WS_E_ENDPOINT_ACTION_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803D0011L))
value WS_E_ENDPOINT_DISCONNECTED (_HRESULT_TYPEDEF_(0x803D0014L))
value WS_E_ENDPOINT_FAILURE (_HRESULT_TYPEDEF_(0x803D000FL))
value WS_E_ENDPOINT_FAULT_RECEIVED (_HRESULT_TYPEDEF_(0x803D0013L))
value WS_E_ENDPOINT_NOT_AVAILABLE (_HRESULT_TYPEDEF_(0x803D000EL))
value WS_E_ENDPOINT_NOT_FOUND (_HRESULT_TYPEDEF_(0x803D000DL))
value WS_E_ENDPOINT_TOO_BUSY (_HRESULT_TYPEDEF_(0x803D0012L))
value WS_E_ENDPOINT_UNREACHABLE (_HRESULT_TYPEDEF_(0x803D0010L))
value WS_E_INVALID_ENDPOINT_URL (_HRESULT_TYPEDEF_(0x803D0020L))
value WS_E_INVALID_FORMAT (_HRESULT_TYPEDEF_(0x803D0000L))
value WS_E_INVALID_OPERATION (_HRESULT_TYPEDEF_(0x803D0003L))
value WS_E_NOT_SUPPORTED (_HRESULT_TYPEDEF_(0x803D0017L))
value WS_E_NO_TRANSLATION_AVAILABLE (_HRESULT_TYPEDEF_(0x803D0009L))
value WS_E_NUMERIC_OVERFLOW (_HRESULT_TYPEDEF_(0x803D0002L))
value WS_E_OBJECT_FAULTED (_HRESULT_TYPEDEF_(0x803D0001L))
value WS_E_OPERATION_ABANDONED (_HRESULT_TYPEDEF_(0x803D0007L))
value WS_E_OPERATION_ABORTED (_HRESULT_TYPEDEF_(0x803D0004L))
value WS_E_OPERATION_TIMED_OUT (_HRESULT_TYPEDEF_(0x803D0006L))
value WS_E_OTHER (_HRESULT_TYPEDEF_(0x803D0021L))
value WS_E_PROXY_ACCESS_DENIED (_HRESULT_TYPEDEF_(0x803D0016L))
value WS_E_PROXY_FAILURE (_HRESULT_TYPEDEF_(0x803D0015L))
value WS_E_PROXY_REQUIRES_BASIC_AUTH (_HRESULT_TYPEDEF_(0x803D0018L))
value WS_E_PROXY_REQUIRES_DIGEST_AUTH (_HRESULT_TYPEDEF_(0x803D0019L))
value WS_E_PROXY_REQUIRES_NEGOTIATE_AUTH (_HRESULT_TYPEDEF_(0x803D001BL))
value WS_E_PROXY_REQUIRES_NTLM_AUTH (_HRESULT_TYPEDEF_(0x803D001AL))
value WS_E_QUOTA_EXCEEDED (_HRESULT_TYPEDEF_(0x803D0008L))
value WS_E_SECURITY_SYSTEM_FAILURE (_HRESULT_TYPEDEF_(0x803D0023L))
value WS_E_SECURITY_TOKEN_EXPIRED (_HRESULT_TYPEDEF_(0x803D0022L))
value WS_E_SECURITY_VERIFICATION_FAILURE (_HRESULT_TYPEDEF_(0x803D000AL))
value WS_E_SERVER_REQUIRES_BASIC_AUTH (_HRESULT_TYPEDEF_(0x803D001CL))
value WS_E_SERVER_REQUIRES_DIGEST_AUTH (_HRESULT_TYPEDEF_(0x803D001DL))
value WS_E_SERVER_REQUIRES_NEGOTIATE_AUTH (_HRESULT_TYPEDEF_(0x803D001FL))
value WS_E_SERVER_REQUIRES_NTLM_AUTH (_HRESULT_TYPEDEF_(0x803D001EL))
value WS_GROUP (0x00020000L)
value WS_HSCROLL (0x00100000L)
value WS_ICONIC (WS_MINIMIZE)
value WS_MAXIMIZE (0x01000000L)
value WS_MAXIMIZEBOX (0x00010000L)
value WS_MINIMIZE (0x20000000L)
value WS_MINIMIZEBOX (0x00020000L)
value WS_OVERLAPPED (0x00000000L)
value WS_OVERLAPPEDWINDOW ((WS_OVERLAPPED | WS_CAPTION | WS_SYSMENU | WS_THICKFRAME | WS_MINIMIZEBOX | WS_MAXIMIZEBOX))
value WS_POPUP (0x80000000L)
value WS_POPUPWINDOW ((WS_POPUP | WS_BORDER | WS_SYSMENU))
value WS_SIZEBOX (WS_THICKFRAME)
value WS_SYSMENU (0x00080000L)
value WS_S_ASYNC (_HRESULT_TYPEDEF_(0x003D0000L))
value WS_S_END (_HRESULT_TYPEDEF_(0x003D0001L))
value WS_TABSTOP (0x00010000L)
value WS_THICKFRAME (0x00040000L)
value WS_TILED (WS_OVERLAPPED)
value WS_TILEDWINDOW (WS_OVERLAPPEDWINDOW)
value WS_VISIBLE (0x10000000L)
value WS_VSCROLL (0x00200000L)
value WTS_CONSOLE_CONNECT (0x1)
value WTS_CONSOLE_DISCONNECT (0x2)
value WTS_REMOTE_CONNECT (0x3)
value WTS_REMOTE_DISCONNECT (0x4)
value WTS_SESSION_CREATE (0xa)
value WTS_SESSION_LOCK (0x7)
value WTS_SESSION_LOGOFF (0x6)
value WTS_SESSION_LOGON (0x5)
value WTS_SESSION_REMOTE_CONTROL (0x9)
value WTS_SESSION_TERMINATE (0xb)
value WTS_SESSION_UNLOCK (0x8)
value WT_EXECUTEDEFAULT (0x00000000)
value WT_EXECUTEDELETEWAIT (0x00000008)
value WT_EXECUTEINIOTHREAD (0x00000001)
value WT_EXECUTEINLONGTHREAD (0x00000010)
value WT_EXECUTEINPERSISTENTIOTHREAD (0x00000040)
value WT_EXECUTEINPERSISTENTTHREAD (0x00000080)
value WT_EXECUTEINTIMERTHREAD (0x00000020)
value WT_EXECUTEINUITHREAD (0x00000002)
value WT_EXECUTEINWAITTHREAD (0x00000004)
value WT_EXECUTELONGFUNCTION (0x00000010)
value WT_EXECUTEONLYONCE (0x00000008)
value WT_TRANSFER_IMPERSONATION (0x00000100)
value WVR_ALIGNBOTTOM (0x0040)
value WVR_ALIGNLEFT (0x0020)
value WVR_ALIGNRIGHT (0x0080)
value WVR_ALIGNTOP (0x0010)
value WVR_HREDRAW (0x0100)
value WVR_REDRAW ((WVR_HREDRAW | WVR_VREDRAW))
value WVR_VALIDRECTS (0x0400)
value WVR_VREDRAW (0x0200)
value XACT_E_ABORTED (_HRESULT_TYPEDEF_(0x8004D019L))
value XACT_E_ABORTING (_HRESULT_TYPEDEF_(0x8004D029L))
value XACT_E_ALREADYINPROGRESS (_HRESULT_TYPEDEF_(0x8004D018L))
value XACT_E_ALREADYOTHERSINGLEPHASE (_HRESULT_TYPEDEF_(0x8004D000L))
value XACT_E_CANTRETAIN (_HRESULT_TYPEDEF_(0x8004D001L))
value XACT_E_CLERKEXISTS (_HRESULT_TYPEDEF_(0x8004D081L))
value XACT_E_CLERKNOTFOUND (_HRESULT_TYPEDEF_(0x8004D080L))
value XACT_E_COMMITFAILED (_HRESULT_TYPEDEF_(0x8004D002L))
value XACT_E_COMMITPREVENTED (_HRESULT_TYPEDEF_(0x8004D003L))
value XACT_E_CONNECTION_DENIED (_HRESULT_TYPEDEF_(0x8004D01DL))
value XACT_E_CONNECTION_DOWN (_HRESULT_TYPEDEF_(0x8004D01CL))
value XACT_E_DEST_TMNOTAVAILABLE (_HRESULT_TYPEDEF_(0x8004D022L))
value XACT_E_FIRST (0x8004D000)
value XACT_E_HEURISTICABORT (_HRESULT_TYPEDEF_(0x8004D004L))
value XACT_E_HEURISTICCOMMIT (_HRESULT_TYPEDEF_(0x8004D005L))
value XACT_E_HEURISTICDAMAGE (_HRESULT_TYPEDEF_(0x8004D006L))
value XACT_E_HEURISTICDANGER (_HRESULT_TYPEDEF_(0x8004D007L))
value XACT_E_INDOUBT (_HRESULT_TYPEDEF_(0x8004D016L))
value XACT_E_INVALIDCOOKIE (_HRESULT_TYPEDEF_(0x8004D015L))
value XACT_E_INVALIDLSN (_HRESULT_TYPEDEF_(0x8004D084L))
value XACT_E_ISOLATIONLEVEL (_HRESULT_TYPEDEF_(0x8004D008L))
value XACT_E_LAST (0x8004D02B)
value XACT_E_LOGFULL (_HRESULT_TYPEDEF_(0x8004D01AL))
value XACT_E_LU_TX_DISABLED (_HRESULT_TYPEDEF_(0x8004D02CL))
value XACT_E_NETWORK_TX_DISABLED (_HRESULT_TYPEDEF_(0x8004D024L))
value XACT_E_NOASYNC (_HRESULT_TYPEDEF_(0x8004D009L))
value XACT_E_NOENLIST (_HRESULT_TYPEDEF_(0x8004D00AL))
value XACT_E_NOIMPORTOBJECT (_HRESULT_TYPEDEF_(0x8004D014L))
value XACT_E_NOISORETAIN (_HRESULT_TYPEDEF_(0x8004D00BL))
value XACT_E_NORESOURCE (_HRESULT_TYPEDEF_(0x8004D00CL))
value XACT_E_NOTCURRENT (_HRESULT_TYPEDEF_(0x8004D00DL))
value XACT_E_NOTIMEOUT (_HRESULT_TYPEDEF_(0x8004D017L))
value XACT_E_NOTRANSACTION (_HRESULT_TYPEDEF_(0x8004D00EL))
value XACT_E_NOTSUPPORTED (_HRESULT_TYPEDEF_(0x8004D00FL))
value XACT_E_PARTNER_NETWORK_TX_DISABLED (_HRESULT_TYPEDEF_(0x8004D025L))
value XACT_E_PULL_COMM_FAILURE (_HRESULT_TYPEDEF_(0x8004D02BL))
value XACT_E_PUSH_COMM_FAILURE (_HRESULT_TYPEDEF_(0x8004D02AL))
value XACT_E_RECOVERYINPROGRESS (_HRESULT_TYPEDEF_(0x8004D082L))
value XACT_E_REENLISTTIMEOUT (_HRESULT_TYPEDEF_(0x8004D01EL))
value XACT_E_REPLAYREQUEST (_HRESULT_TYPEDEF_(0x8004D085L))
value XACT_E_TIP_CONNECT_FAILED (_HRESULT_TYPEDEF_(0x8004D01FL))
value XACT_E_TIP_DISABLED (_HRESULT_TYPEDEF_(0x8004D023L))
value XACT_E_TIP_PROTOCOL_ERROR (_HRESULT_TYPEDEF_(0x8004D020L))
value XACT_E_TIP_PULL_FAILED (_HRESULT_TYPEDEF_(0x8004D021L))
value XACT_E_TMNOTAVAILABLE (_HRESULT_TYPEDEF_(0x8004D01BL))
value XACT_E_TRANSACTIONCLOSED (_HRESULT_TYPEDEF_(0x8004D083L))
value XACT_E_UNABLE_TO_LOAD_DTC_PROXY (_HRESULT_TYPEDEF_(0x8004D028L))
value XACT_E_UNABLE_TO_READ_DTC_CONFIG (_HRESULT_TYPEDEF_(0x8004D027L))
value XACT_E_UNKNOWNRMGRID (_HRESULT_TYPEDEF_(0x8004D010L))
value XACT_E_WRONGSTATE (_HRESULT_TYPEDEF_(0x8004D011L))
value XACT_E_WRONGUOW (_HRESULT_TYPEDEF_(0x8004D012L))
value XACT_E_XA_TX_DISABLED (_HRESULT_TYPEDEF_(0x8004D026L))
value XACT_E_XTIONEXISTS (_HRESULT_TYPEDEF_(0x8004D013L))
value XACT_S_ABORTING (_HRESULT_TYPEDEF_(0x0004D008L))
value XACT_S_ALLNORETAIN (_HRESULT_TYPEDEF_(0x0004D007L))
value XACT_S_ASYNC (_HRESULT_TYPEDEF_(0x0004D000L))
value XACT_S_DEFECT (_HRESULT_TYPEDEF_(0x0004D001L))
value XACT_S_FIRST (0x0004D000)
value XACT_S_LAST (0x0004D010)
value XACT_S_LASTRESOURCEMANAGER (_HRESULT_TYPEDEF_(0x0004D010L))
value XACT_S_LOCALLY_OK (_HRESULT_TYPEDEF_(0x0004D00AL))
value XACT_S_MADECHANGESCONTENT (_HRESULT_TYPEDEF_(0x0004D005L))
value XACT_S_MADECHANGESINFORM (_HRESULT_TYPEDEF_(0x0004D006L))
value XACT_S_OKINFORM (_HRESULT_TYPEDEF_(0x0004D004L))
value XACT_S_READONLY (_HRESULT_TYPEDEF_(0x0004D002L))
value XACT_S_SINGLEPHASE (_HRESULT_TYPEDEF_(0x0004D009L))
value XACT_S_SOMENORETAIN (_HRESULT_TYPEDEF_(0x0004D003L))
value XCLASS_BOOL (0x1000)
value XCLASS_DATA (0x2000)
value XCLASS_FLAGS (0x4000)
value XCLASS_MASK (0xFC00)
value XCLASS_NOTIFICATION (0x8000)
value XENROLL_E_CANNOT_ADD_ROOT_CERT (_HRESULT_TYPEDEF_(0x80095001L))
value XENROLL_E_KEYSPEC_SMIME_MISMATCH (_HRESULT_TYPEDEF_(0x80095005L))
value XENROLL_E_KEY_NOT_EXPORTABLE (_HRESULT_TYPEDEF_(0x80095000L))
value XENROLL_E_RESPONSE_KA_HASH_MISMATCH (_HRESULT_TYPEDEF_(0x80095004L))
value XENROLL_E_RESPONSE_KA_HASH_NOT_FOUND (_HRESULT_TYPEDEF_(0x80095002L))
value XENROLL_E_RESPONSE_UNEXPECTED_KA_HASH (_HRESULT_TYPEDEF_(0x80095003L))
value XSTATE_ALIGN_BIT ((1))
value XSTATE_AMX_TILE_CONFIG ((17))
value XSTATE_AMX_TILE_DATA ((18))
value XSTATE_AVX ((XSTATE_GSSE))
value XSTATE_CET_S ((12))
value XSTATE_CET_U ((11))
value XSTATE_COMPACTION_ENABLE ((63))
value XSTATE_CONTROLFLAG_VALID_MASK ((XSTATE_CONTROLFLAG_XSAVEOPT_MASK | XSTATE_CONTROLFLAG_XSAVEC_MASK | XSTATE_CONTROLFLAG_XFD_MASK))
value XSTATE_CONTROLFLAG_XFD_MASK ((4))
value XSTATE_CONTROLFLAG_XSAVEC_MASK ((2))
value XSTATE_CONTROLFLAG_XSAVEOPT_MASK ((1))
value XSTATE_GSSE ((2))
value XSTATE_IPT ((8))
value XSTATE_LEGACY_FLOATING_POINT ((0))
value XSTATE_LEGACY_SSE ((1))
value XSTATE_LWP ((62))
value XSTATE_MASK_ALLOWED ((XSTATE_MASK_LEGACY | XSTATE_MASK_AVX | XSTATE_MASK_MPX | XSTATE_MASK_AVX512 | XSTATE_MASK_IPT | XSTATE_MASK_PASID | XSTATE_MASK_CET_U | XSTATE_MASK_AMX_TILE_CONFIG | XSTATE_MASK_AMX_TILE_DATA | XSTATE_MASK_LWP))
value XSTATE_MASK_AVX ((XSTATE_MASK_GSSE))
value XSTATE_MASK_LARGE_FEATURES ((XSTATE_MASK_AMX_TILE_DATA))
value XSTATE_MASK_LEGACY ((XSTATE_MASK_LEGACY_FLOATING_POINT | XSTATE_MASK_LEGACY_SSE))
value XSTATE_MASK_USER_VISIBLE_SUPERVISOR ((XSTATE_MASK_CET_U))
value XSTATE_MPX_BNDCSR ((4))
value XSTATE_MPX_BNDREGS ((3))
value XSTATE_PASID ((10))
value XSTATE_XFD_BIT ((2))
value XST_ADVACKRCVD (13)
value XST_ADVDATAACKRCVD (16)
value XST_ADVDATASENT (15)
value XST_ADVSENT (11)
value XST_CONNECTED (2)
value XST_DATARCVD (6)
value XST_EXECACKRCVD (10)
value XST_EXECSENT (9)
value XST_INCOMPLETE (1)
value XST_NULL (0)
value XST_POKEACKRCVD (8)
value XST_POKESENT (7)
value XST_REQSENT (5)
value XST_UNADVACKRCVD (14)
value XST_UNADVSENT (12)
value XTYPF_ACKREQ (0x0008)
value XTYPF_NOBLOCK (0x0002)
value XTYPF_NODATA (0x0004)
value XTYP_ADVDATA ((0x0010 | XCLASS_FLAGS ))
value XTYP_ADVREQ ((0x0020 | XCLASS_DATA | XTYPF_NOBLOCK ))
value XTYP_ADVSTART ((0x0030 | XCLASS_BOOL ))
value XTYP_ADVSTOP ((0x0040 | XCLASS_NOTIFICATION))
value XTYP_CONNECT ((0x0060 | XCLASS_BOOL | XTYPF_NOBLOCK))
value XTYP_CONNECT_CONFIRM ((0x0070 | XCLASS_NOTIFICATION | XTYPF_NOBLOCK))
value XTYP_DISCONNECT ((0x00C0 | XCLASS_NOTIFICATION | XTYPF_NOBLOCK))
value XTYP_ERROR ((0x0000 | XCLASS_NOTIFICATION | XTYPF_NOBLOCK ))
value XTYP_EXECUTE ((0x0050 | XCLASS_FLAGS ))
value XTYP_MASK (0x00F0)
value XTYP_MONITOR ((0x00F0 | XCLASS_NOTIFICATION | XTYPF_NOBLOCK))
value XTYP_POKE ((0x0090 | XCLASS_FLAGS ))
value XTYP_REGISTER ((0x00A0 | XCLASS_NOTIFICATION | XTYPF_NOBLOCK))
value XTYP_REQUEST ((0x00B0 | XCLASS_DATA ))
value XTYP_SHIFT (4)
value XTYP_UNREGISTER ((0x00D0 | XCLASS_NOTIFICATION | XTYPF_NOBLOCK))
value XTYP_WILDCONNECT ((0x00E0 | XCLASS_DATA | XTYPF_NOBLOCK))
value XTYP_XACT_COMPLETE ((0x0080 | XCLASS_NOTIFICATION ))
value ZAWPROXYAPI (DECLSPEC_IMPORT)
value ZERO_PADDING (3)
value _ACRTIMP_ALT (_ACRTIMP)
value _ALPHA ((0x0100 | _UPPER | _LOWER))
value _ARGMAX (100)
value _ARM_WINAPI_PARTITION_DESKTOP_SDK_AVAILABLE (1)
value _ASSEMBLY_DLL_REDIRECTION_DETAILED_INFORMATION (_ASSEMBLY_FILE_DETAILED_INFORMATION)
value _BLANK (0x40)
value _CALL_REPORTFAULT (0x2)
value _CONTROL (0x20)
value _CRT_BUILD_DESKTOP_APP (1)
value _CRT_FUNCTIONS_REQUIRED (1)
value _CRT_INTERNAL_NONSTDC_NAMES (1)
value _CRT_INT_MAX (2147483647)
value _CRT_PACKING (8)
value _CRT_SECURE_CPP_OVERLOAD_SECURE_NAMES (1)
value _CRT_SECURE_CPP_OVERLOAD_SECURE_NAMES_MEMORY (0)
value _CRT_SECURE_CPP_OVERLOAD_STANDARD_NAMES (0)
value _CRT_SECURE_CPP_OVERLOAD_STANDARD_NAMES_COUNT (0)
value _CRT_SECURE_CPP_OVERLOAD_STANDARD_NAMES_MEMORY (0)
value _CRT_USE_CONFORMING_ANNEX_K_TIME (0)
value _CVTBUFSIZE ((309 + 40))
value _DIGIT (0x04)
value _HAS_EXCEPTIONS (1)
value _HAS_NODISCARD (0)
value _HEX (0x80)
value _INTEGRAL_MAX_BITS (64)
value _IOB_ENTRIES (3)
value _IOFBF (0x0000)
value _IOLBF (0x0040)
value _IONBF (0x0004)
value _LEADBYTE (0x8000)
value _LOWER (0x02)
value _MAX_DIR (256)
value _MAX_DRIVE (3)
value _MAX_ENV (32767)
value _MAX_EXT (256)
value _MAX_FNAME (256)
value _MAX_PATH (260)
value _MM_HINT_NTA (0)
value _MSC_BUILD (1)
value _MSC_EXTENSIONS (1)
value _MSC_FULL_VER (192000000)
value _MSC_VER (1920)
value _MSVC_EXECUTION_CHARACTER_SET (65001)
value _NFILE (_NSTREAM_)
value _NLSCMPERROR (_CRT_INT_MAX)
value _NSTREAM_ (512)
value _OUT_TO_DEFAULT (0)
value _OUT_TO_MSGBOX (2)
value _OUT_TO_STDERR (1)
value _O_APPEND (0x0008)
value _O_BINARY (0x8000)
value _O_CREAT (0x0100)
value _O_EXCL (0x0400)
value _O_NOINHERIT (0x0080)
value _O_OBTAIN_DIR (0x2000)
value _O_RANDOM (0x0010)
value _O_RAW (_O_BINARY)
value _O_RDONLY (0x0000)
value _O_RDWR (0x0002)
value _O_SEQUENTIAL (0x0020)
value _O_SHORT_LIVED (0x1000)
value _O_TEMPORARY (0x0040)
value _O_TEXT (0x4000)
value _O_TRUNC (0x0200)
value _O_WRONLY (0x0001)
value _O_WTEXT (0x10000)
value _PUNCT (0x10)
value _REPORT_ERRMODE (3)
value _RPC_HTTP_TRANSPORT_CREDENTIALS (_RPC_HTTP_TRANSPORT_CREDENTIALS_A)
value _SAL_VERSION (20)
value _SECURECRT_FILL_BUFFER_PATTERN (0xFE)
value _SEC_WINNT_AUTH_IDENTITY (_SEC_WINNT_AUTH_IDENTITY_A)
value _SPACE (0x08)
value _SS_MAXSIZE (128)
value _STRALIGN_USE_SECURE_CRT (1)
value _SYS_OPEN (20)
value _S_IEXEC (0x0040)
value _S_IFCHR (0x2000)
value _S_IFDIR (0x4000)
value _S_IFIFO (0x1000)
value _S_IFMT (0xF000)
value _S_IFREG (0x8000)
value _S_IREAD (0x0100)
value _S_IWRITE (0x0080)
value _TMP_MAX_S (TMP_MAX)
value _UCRT_DISABLED_WARNINGS (4324 _UCRT_DISABLED_WARNING_4412 4514 4574 4710 4793 4820 4995 4996 28719 28726 28727 _UCRT_EXTRA_DISABLED_WARNINGS)
value _UPPER (0x01)
value _USE_ATTRIBUTES_FOR_SAL (0)
value _USE_DECLSPECS_FOR_SAL (0)
value _VCRT_COMPILER_PREPROCESSOR (1)
value _VCRUNTIME_DISABLED_WARNINGS (_VCRUNTIME_DISABLED_WARNING_4339 _VCRUNTIME_DISABLED_WARNING_4412 4514 4820 _VCRUNTIME_EXTRA_DISABLED_WARNINGS)
value _WRITE_ABORT_MSG (0x1)
value __ATOMIC_ACQUIRE (2)
value __ATOMIC_ACQ_REL (4)
value __ATOMIC_CONSUME (1)
value __ATOMIC_RELAXED (0)
value __ATOMIC_RELEASE (3)
value __ATOMIC_SEQ_CST (5)
value __BIGGEST_ALIGNMENT__ (16)
value __BITINT_MAXWIDTH__ (128)
value __BOOL_WIDTH__ (8)
value __BYTE_ORDER__ (__ORDER_LITTLE_ENDIAN__)
value __CHAR_BIT__ (8)
value __CLANG_ATOMIC_BOOL_LOCK_FREE (2)
value __CLANG_ATOMIC_CHAR_LOCK_FREE (2)
value __CLANG_ATOMIC_INT_LOCK_FREE (2)
value __CLANG_ATOMIC_LLONG_LOCK_FREE (2)
value __CLANG_ATOMIC_LONG_LOCK_FREE (2)
value __CLANG_ATOMIC_POINTER_LOCK_FREE (2)
value __CLANG_ATOMIC_SHORT_LOCK_FREE (2)
value __CLANG_ATOMIC_WCHAR_T_LOCK_FREE (2)
value __CONSTANT_CFSTRINGS__ (1)
value __CRTDECL (__CLRCALL_PURE_OR_CDECL)
value __DBL_DECIMAL_DIG__ (17)
value __DBL_DIG__ (15)
value __DBL_HAS_DENORM__ (1)
value __DBL_HAS_INFINITY__ (1)
value __DBL_HAS_QUIET_NAN__ (1)
value __DBL_MANT_DIG__ (53)
value __DBL_MAX_EXP__ (1024)
value __DBL_MIN_EXP__ ((-1021))
value __DECIMAL_DIG__ (__LDBL_DECIMAL_DIG__)
value __FILEW__ (_CRT_WIDE(__FILE__))
value __FINITE_MATH_ONLY__ (0)
value __FLT_DECIMAL_DIG__ (9)
value __FLT_DIG__ (6)
value __FLT_HAS_DENORM__ (1)
value __FLT_HAS_INFINITY__ (1)
value __FLT_HAS_QUIET_NAN__ (1)
value __FLT_MANT_DIG__ (24)
value __FLT_MAX_EXP__ (128)
value __FLT_MIN_EXP__ ((-125))
value __FLT_RADIX__ (2)
value __FUNCTIONW__ (_CRT_WIDE(__FUNCTION__))
value __FXSR__ (1)
value __GCC_ASM_FLAG_OUTPUTS__ (1)
value __GOT_SECURE_LIB__ (__STDC_SECURE_LIB__)
value __INTMAX_C_SUFFIX__ (LL)
value __INTMAX_MAX__ (9223372036854775807LL)
value __INTMAX_WIDTH__ (64)
value __INTPTR_MAX__ (9223372036854775807LL)
value __INTPTR_WIDTH__ (64)
value __INT_MAX__ (2147483647)
value __INT_WIDTH__ (32)
value __LDBL_DECIMAL_DIG__ (17)
value __LDBL_DIG__ (15)
value __LDBL_HAS_DENORM__ (1)
value __LDBL_HAS_INFINITY__ (1)
value __LDBL_HAS_QUIET_NAN__ (1)
value __LDBL_MANT_DIG__ (53)
value __LDBL_MAX_EXP__ (1024)
value __LDBL_MIN_EXP__ ((-1021))
value __LITTLE_ENDIAN__ (1)
value __LLONG_WIDTH__ (64)
value __LONG_LONG_MAX__ (9223372036854775807LL)
value __LONG_MAX__ (2147483647)
value __LONG_WIDTH__ (32)
value __MMX__ (1)
value __NO_INLINE__ (1)
value __NO_MATH_INLINES (1)
value __OBJC_BOOL_IS_BOOL (0)
value __OPENCL_MEMORY_SCOPE_ALL_SVM_DEVICES (3)
value __OPENCL_MEMORY_SCOPE_DEVICE (2)
value __OPENCL_MEMORY_SCOPE_SUB_GROUP (4)
value __OPENCL_MEMORY_SCOPE_WORK_GROUP (1)
value __OPENCL_MEMORY_SCOPE_WORK_ITEM (0)
value __ORDER_BIG_ENDIAN__ (4321)
value __ORDER_LITTLE_ENDIAN__ (1234)
value __ORDER_PDP_ENDIAN__ (3412)
value __PIC__ (2)
value __POINTER_WIDTH__ (64)
value __PRAGMA_REDEFINE_EXTNAME (1)
value __PTRDIFF_MAX__ (9223372036854775807LL)
value __PTRDIFF_WIDTH__ (64)
value __REQUIRED_RPCNDR_H_VERSION__ (501)
value __REQUIRED_RPCSAL_H_VERSION__ (100)
value __RPCNDR_H_VERSION__ (( 501 ))
value __RPCSAL_H_VERSION__ (( 100 ))
value __SAL_H_FULL_VER (140050727)
value __SAL_H_VERSION (180000000)
value __SCHAR_MAX__ (127)
value __SEG_FS (1)
value __SEG_GS (1)
value __SHRT_MAX__ (32767)
value __SHRT_WIDTH__ (16)
value __SIG_ATOMIC_MAX__ (2147483647)
value __SIG_ATOMIC_WIDTH__ (32)
value __SIZEOF_DOUBLE__ (8)
value __SIZEOF_FLOAT__ (4)
value __SIZEOF_INT__ (4)
value __SIZEOF_LONG_DOUBLE__ (8)
value __SIZEOF_LONG_LONG__ (8)
value __SIZEOF_LONG__ (4)
value __SIZEOF_POINTER__ (8)
value __SIZEOF_PTRDIFF_T__ (8)
value __SIZEOF_SHORT__ (2)
value __SIZEOF_SIZE_T__ (8)
value __SIZEOF_WCHAR_T__ (2)
value __SIZEOF_WINT_T__ (2)
value __SIZE_MAX__ (18446744073709551615ULL)
value __SIZE_WIDTH__ (64)
value __SPECSTRINGS_STRICT_LEVEL (1)
value __SSE_MATH__ (1)
value __SSE__ (1)
value __STDC_HOSTED__ (1)
value __STDC_NO_THREADS__ (1)
value __STDC_SECURE_LIB__ (200411)
value __STDC_VERSION__ (201710)
value __STDC_WANT_SECURE_LIB__ (1)
value __UINTMAX_C_SUFFIX__ (ULL)
value __UINTMAX_MAX__ (18446744073709551615ULL)
value __UINTMAX_WIDTH__ (64)
value __UINTPTR_MAX__ (18446744073709551615ULL)
value __UINTPTR_WIDTH__ (64)
value __WCHAR_MAX__ (65535)
value __WCHAR_UNSIGNED__ (1)
value __WCHAR_WIDTH__ (16)
value __WINT_MAX__ (65535)
value __WINT_UNSIGNED__ (1)
value __WINT_WIDTH__ (16)

