
value EAGAIN (536870918)
value SOCK_STREAM (1)

value SOL_SOCKET (65535)
value SO_REUSEADDR (4)
value SO_RCVTIMEO (4102)

value AF_INET (2)
value AF_UNIX (1)

value AI_PASSIVE (1)
value AI_CANONNAME (2)
value AI_NUMERICHOST (4)

value POLLIN (768)
value POLLOUT (16)
value POLLERR (1)
value POLLHUP (2)

value WSAENOBUFS (10055)
value FIONBIO (2148034174)