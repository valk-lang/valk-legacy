
value ABE_BOTTOM (3)
value ABE_LEFT (0)
value ABE_RIGHT (2)
value ABE_TOP (1)
value ABORTDOC (2)
value ABSOLUTE (1)
value ACCESS_MAX_LEVEL (4)
value ACCESS_OBJECT_GUID (0)
value ACCESS_PROPERTY_GUID (2)
value ACCESS_PROPERTY_SET_GUID (1)
value ACTIVATIONCONTEXTINFOCLASS (ACTIVATION_CONTEXT_INFO_CLASS)
value ACTIVATION_CONTEXT_BASIC_INFORMATION_DEFINED (1)
value ADDR_ANY (INADDR_ANY)
value AD_CLOCKWISE (2)
value AD_COUNTERCLOCKWISE (1)
value AF_APPLETALK (16)
value AF_ATM (22)
value AF_BAN (21)
value AF_BTH (32)
value AF_CCITT (10)
value AF_CHAOS (5)
value AF_CLUSTER (24)
value AF_DATAKIT (9)
value AF_DLI (13)
value AF_ECMA (8)
value AF_FIREFOX (19)
value AF_HYLINK (15)
value AF_HYPERV (34)
value AF_ICLFXBM (31)
value AF_IMPLINK (3)
value AF_INET (2)
value AF_IPX (AF_NS)
value AF_IRDA (26)
value AF_ISO (7)
value AF_LAT (14)
value AF_LINK (33)
value AF_MAX (35)
value AF_NETBIOS (17)
value AF_NETDES (28)
value AF_NS (6)
value AF_OSI (AF_ISO)
value AF_PUP (4)
value AF_SNA (11)
value AF_TCNMESSAGE (30)
value AF_TCNPROCESS (29)
value AF_UNIX (1)
value AF_UNSPEC (0)
value AF_VOICEVIEW (18)
value ALERT_SYSTEM_CRITICAL (5)
value ALERT_SYSTEM_ERROR (3)
value ALERT_SYSTEM_INFORMATIONAL (1)
value ALERT_SYSTEM_QUERY (4)
value ALERT_SYSTEM_WARNING (2)
value ALG_SID_AES (17)
value ALG_SID_AGREED_KEY_ANY (3)
value ALG_SID_CAST (6)
value ALG_SID_CYLINK_MEK (12)
value ALG_SID_DES (1)
value ALG_SID_DESX (4)
value ALG_SID_DH_EPHEM (2)
value ALG_SID_DH_SANDF (1)
value ALG_SID_DSS_ANY (0)
value ALG_SID_DSS_DMS (2)
value ALG_SID_DSS_PKCS (1)
value ALG_SID_ECDH (5)
value ALG_SID_ECDH_EPHEM (6)
value ALG_SID_ECDSA (3)
value ALG_SID_ECMQV (1)
value ALG_SID_EXAMPLE (80)
value ALG_SID_HASH_REPLACE_OWF (11)
value ALG_SID_HMAC (9)
value ALG_SID_IDEA (5)
value ALG_SID_KEA (4)
value ALG_SID_MAC (5)
value ALG_SID_RIPEMD (6)
value ALG_SID_RSA_ANY (0)
value ALG_SID_RSA_ENTRUST (3)
value ALG_SID_RSA_MSATWORK (2)
value ALG_SID_RSA_PGP (4)
value ALG_SID_RSA_PKCS (1)
value ALG_SID_SCHANNEL_ENC_KEY (7)
value ALG_SID_SCHANNEL_MAC_KEY (3)
value ALG_SID_SCHANNEL_MASTER_HASH (2)
value ALG_SID_SEAL (2)
value ALG_SID_SHA (4)
value ALG_SID_SKIPJACK (10)
value ALG_SID_TEK (11)
value ALTERNATE (1)
value ANSI_CHARSET (0)
value ANSI_FIXED_FONT (11)
value ANSI_VAR_FONT (12)
value ANTIALIASED_QUALITY (4)
value ANYSIZE_ARRAY (1)
value APC_LEVEL (1)
value APIENTRY (WINAPI)
value APPCOMMAND_BASS_BOOST (20)
value APPCOMMAND_BASS_DOWN (19)
value APPCOMMAND_BASS_UP (21)
value APPCOMMAND_BROWSER_BACKWARD (1)
value APPCOMMAND_BROWSER_FAVORITES (6)
value APPCOMMAND_BROWSER_FORWARD (2)
value APPCOMMAND_BROWSER_HOME (7)
value APPCOMMAND_BROWSER_REFRESH (3)
value APPCOMMAND_BROWSER_SEARCH (5)
value APPCOMMAND_BROWSER_STOP (4)
value APPCOMMAND_CLOSE (31)
value APPCOMMAND_COPY (36)
value APPCOMMAND_CORRECTION_LIST (45)
value APPCOMMAND_CUT (37)
value APPCOMMAND_DELETE (53)
value APPCOMMAND_DICTATE_OR_COMMAND_CONTROL_TOGGLE (43)
value APPCOMMAND_FIND (28)
value APPCOMMAND_FORWARD_MAIL (40)
value APPCOMMAND_HELP (27)
value APPCOMMAND_LAUNCH_MAIL (15)
value APPCOMMAND_LAUNCH_MEDIA_SELECT (16)
value APPCOMMAND_MEDIA_CHANNEL_DOWN (52)
value APPCOMMAND_MEDIA_CHANNEL_UP (51)
value APPCOMMAND_MEDIA_FAST_FORWARD (49)
value APPCOMMAND_MEDIA_NEXTTRACK (11)
value APPCOMMAND_MEDIA_PAUSE (47)
value APPCOMMAND_MEDIA_PLAY (46)
value APPCOMMAND_MEDIA_PLAY_PAUSE (14)
value APPCOMMAND_MEDIA_PREVIOUSTRACK (12)
value APPCOMMAND_MEDIA_RECORD (48)
value APPCOMMAND_MEDIA_REWIND (50)
value APPCOMMAND_MEDIA_STOP (13)
value APPCOMMAND_MICROPHONE_VOLUME_DOWN (25)
value APPCOMMAND_MICROPHONE_VOLUME_MUTE (24)
value APPCOMMAND_MICROPHONE_VOLUME_UP (26)
value APPCOMMAND_MIC_ON_OFF_TOGGLE (44)
value APPCOMMAND_NEW (29)
value APPCOMMAND_OPEN (30)
value APPCOMMAND_PASTE (38)
value APPCOMMAND_PRINT (33)
value APPCOMMAND_REDO (35)
value APPCOMMAND_REPLY_TO_MAIL (39)
value APPCOMMAND_SAVE (32)
value APPCOMMAND_SEND_MAIL (41)
value APPCOMMAND_SPELL_CHECK (42)
value APPCOMMAND_TREBLE_DOWN (22)
value APPCOMMAND_TREBLE_UP (23)
value APPCOMMAND_UNDO (34)
value APPCOMMAND_VOLUME_DOWN (9)
value APPCOMMAND_VOLUME_MUTE (8)
value APPCOMMAND_VOLUME_UP (10)
value APPMODEL_ERROR_DYNAMIC_PROPERTY_INVALID (15705L)
value APPMODEL_ERROR_DYNAMIC_PROPERTY_READ_FAILED (15704L)
value APPMODEL_ERROR_NO_APPLICATION (15703L)
value APPMODEL_ERROR_NO_MUTABLE_DIRECTORY (15707L)
value APPMODEL_ERROR_NO_PACKAGE (15700L)
value APPMODEL_ERROR_PACKAGE_IDENTITY_CORRUPT (15702L)
value APPMODEL_ERROR_PACKAGE_NOT_AVAILABLE (15706L)
value APPMODEL_ERROR_PACKAGE_RUNTIME_CORRUPT (15701L)
value APP_LOCAL_DEVICE_ID_SIZE (32)
value ARABIC_CHARSET (178)
value ARM_CACHE_ALIGNMENT_SIZE (128)
value ASPECTX (40)
value ASPECTXY (44)
value ASPECTY (42)
value ASSEMBLY_DLL_REDIRECTION_DETAILED_INFORMATION (ASSEMBLY_FILE_DETAILED_INFORMATION)
value AT_KEYEXCHANGE (1)
value AT_SIGNATURE (2)
value AUTHTYPE_CLIENT (1)
value AUTHTYPE_SERVER (2)
value AUXCAPS_AUXIN (2)
value AUXCAPS_CDAUDIO (1)
value BALTIC_CHARSET (186)
value BANDINFO (24)
value BASE_PROTOCOL (1)
value BCRYPTBUFFER_VERSION (0)
value BCRYPT_AUTHENTICATED_CIPHER_MODE_INFO_VERSION (1)
value BCRYPT_OBJECT_ALIGNMENT (16)
value BEGIN_PATH (4096)
value BINDF_DONTPUTINCACHE (BINDF_NOWRITECACHE)
value BINDF_DONTUSECACHE (BINDF_GETNEWESTVERSION)
value BINDF_NOCOPYDATA (BINDF_PULLDATA)
value BITSPIXEL (12)
value BI_BITFIELDS (3L)
value BI_JPEG (4L)
value BI_PNG (5L)
value BI_RGB (0cL)
value BKMODE_LAST (2)
value BLACKONWHITE (1)
value BLACK_BRUSH (4)
value BLACK_PEN (7)
value BLTALIGNMENT (119)
value BN_CLICKED (0)
value BN_DBLCLK (BN_DOUBLECLICKED)
value BN_DISABLE (4)
value BN_DOUBLECLICKED (5)
value BN_HILITE (2)
value BN_KILLFOCUS (7)
value BN_PAINT (1)
value BN_PUSHED (BN_HILITE)
value BN_SETFOCUS (6)
value BN_UNHILITE (3)
value BN_UNPUSHED (BN_UNHILITE)
value BS_DIBPATTERN (5)
value BS_DIBPATTERNPT (6)
value BS_HATCHED (2)
value BS_HOLLOW (BS_NULL)
value BS_INDEXED (4)
value BS_MONOPATTERN (9)
value BS_NULL (1)
value BS_PATTERN (3)
value BS_RIGHTBUTTON (BS_LEFTTEXT)
value BS_SOLID (0)
value BUFSIZ (512)
value CALERT_SYSTEM (6)
value CALINFO_ENUMPROC (CALINFO_ENUMPROCA)
value CALINFO_ENUMPROCEX (CALINFO_ENUMPROCEXA)
value CAL_GREGORIAN (1)
value CAL_GREGORIAN_ARABIC (10)
value CAL_GREGORIAN_ME_FRENCH (9)
value CAL_GREGORIAN_US (2)
value CAL_GREGORIAN_XLIT_ENGLISH (11)
value CAL_GREGORIAN_XLIT_FRENCH (12)
value CAL_HEBREW (8)
value CAL_HIJRI (6)
value CAL_JAPAN (3)
value CAL_KOREA (5)
value CAL_NOUSEROVERRIDE (LOCALE_NOUSEROVERRIDE)
value CAL_PERSIAN (22)
value CAL_RETURN_GENITIVE_NAMES (LOCALE_RETURN_GENITIVE_NAMES)
value CAL_RETURN_NUMBER (LOCALE_RETURN_NUMBER)
value CAL_TAIWAN (4)
value CAL_THAI (7)
value CAL_UMALQURA (23)
value CAL_USE_CP_ACP (LOCALE_USE_CP_ACP)
value CAP_ATAPI_ID_CMD (2)
value CAP_ATA_ID_CMD (1)
value CAP_SMART_CMD (4)
value CBN_CLOSEUP (8)
value CBN_DBLCLK (2)
value CBN_DROPDOWN (7)
value CBN_EDITCHANGE (5)
value CBN_EDITUPDATE (6)
value CBN_KILLFOCUS (4)
value CBN_SELCHANGE (1)
value CBN_SELENDCANCEL (10)
value CBN_SELENDOK (9)
value CBN_SETFOCUS (3)
value CB_OKAY (0)
value CCHDEVICENAME (32)
value CCHFORMNAME (32)
value CCHILDREN_SCROLLBAR (5)
value CCHILDREN_TITLEBAR (5)
value CCH_MAX_PROPSTG_NAME (31)
value CC_CHORD (4)
value CC_CIRCLES (1)
value CC_ELLIPSES (8)
value CC_INTERIORS (128)
value CC_NONE (0)
value CC_PIE (2)
value CC_ROUNDRECT (256)
value CC_STYLED (32)
value CC_WIDE (16)
value CC_WIDESTYLED (64)
value CDB_SIZE (16)
value CD_LBSELADD (2)
value CD_LBSELCHANGE (0)
value CD_LBSELSUB (1)
value CERT_ACCESS_STATE_PROP_ID (14)
value CERT_AIA_URL_RETRIEVED_PROP_ID (67)
value CERT_ALT_NAME_DIRECTORY_NAME (5)
value CERT_ALT_NAME_DNS_NAME (3)
value CERT_ALT_NAME_EDI_PARTY_NAME (6)
value CERT_ALT_NAME_ENTRY_ERR_INDEX_SHIFT (16)
value CERT_ALT_NAME_IP_ADDRESS (8)
value CERT_ALT_NAME_OTHER_NAME (1)
value CERT_ALT_NAME_REGISTERED_ID (9)
value CERT_ALT_NAME_URL (7)
value CERT_ALT_NAME_VALUE_ERR_INDEX_SHIFT (0)
value CERT_ARCHIVED_KEY_HASH_PROP_ID (65)
value CERT_ARCHIVED_PROP_ID (19)
value CERT_AUTHORITY_INFO_ACCESS_PROP_ID (68)
value CERT_AUTH_ROOT_AUTO_UPDATE_LOCAL_MACHINE_REGPATH (CERT_AUTO_UPDATE_LOCAL_MACHINE_REGPATH)
value CERT_AUTH_ROOT_AUTO_UPDATE_ROOT_DIR_URL_VALUE_NAME (CERT_AUTO_UPDATE_ROOT_DIR_URL_VALUE_NAME)
value CERT_AUTO_ENROLL_PROP_ID (21)
value CERT_AUTO_ENROLL_RETRY_PROP_ID (66)
value CERT_BACKED_UP_PROP_ID (69)
value CERT_BIOMETRIC_OID_DATA_CHOICE (2)
value CERT_BIOMETRIC_PICTURE_TYPE (0)
value CERT_BIOMETRIC_PREDEFINED_DATA_CHOICE (1)
value CERT_BIOMETRIC_SIGNATURE_TYPE (1)
value CERT_BUNDLE_CERTIFICATE (0)
value CERT_BUNDLE_CRL (1)
value CERT_CA_DISABLE_CRL_PROP_ID (82)
value CERT_CA_OCSP_AUTHORITY_INFO_ACCESS_PROP_ID (81)
value CERT_CEP_PROP_ID (87)
value CERT_CHAIN_AUTO_CURRENT_USER (1)
value CERT_CHAIN_AUTO_HPKP_RULE_INFO (8)
value CERT_CHAIN_AUTO_IMPERSONATED (3)
value CERT_CHAIN_AUTO_LOCAL_MACHINE (2)
value CERT_CHAIN_AUTO_NETWORK_INFO (6)
value CERT_CHAIN_AUTO_PINRULE_INFO (5)
value CERT_CHAIN_AUTO_PROCESS_INFO (4)
value CERT_CHAIN_AUTO_SERIAL_LOCAL_MACHINE (7)
value CERT_CHAIN_CRL_VALIDITY_EXT_PERIOD_HOURS_DEFAULT (12)
value CERT_CHAIN_FIND_BY_ISSUER (1)
value CERT_CHAIN_MAX_AIA_URL_COUNT_IN_CERT_DEFAULT (5)
value CERT_CHAIN_MAX_AIA_URL_RETRIEVAL_BYTE_COUNT_DEFAULT (100000)
value CERT_CHAIN_MAX_AIA_URL_RETRIEVAL_CERT_COUNT_DEFAULT (10)
value CERT_CHAIN_MAX_AIA_URL_RETRIEVAL_COUNT_PER_CHAIN_DEFAULT (3)
value CERT_CHAIN_MAX_SSL_TIME_UPDATED_EVENT_COUNT_DEFAULT (5)
value CERT_CHAIN_MIN_RSA_PUB_KEY_BIT_LENGTH_DEFAULT (1023)
value CERT_CHAIN_POLICY_SSL_KEY_PIN_MISMATCH_WARNING (2)
value CERT_CHAIN_POLICY_SSL_KEY_PIN_MITM_WARNING (1)
value CERT_CHAIN_POLICY_SSL_KEY_PIN_SUCCESS (0)
value CERT_CLR_DELETE_KEY_PROP_ID (125)
value CERT_COMPARE_ANY (0)
value CERT_COMPARE_ATTR (3)
value CERT_COMPARE_CERT_ID (16)
value CERT_COMPARE_CROSS_CERT_DIST_POINTS (17)
value CERT_COMPARE_CTL_USAGE (CERT_COMPARE_ENHKEY_USAGE)
value CERT_COMPARE_ENHKEY_USAGE (10)
value CERT_COMPARE_EXISTING (13)
value CERT_COMPARE_HASH (CERT_COMPARE_SHA1_HASH)
value CERT_COMPARE_HASH_STR (20)
value CERT_COMPARE_HAS_PRIVATE_KEY (21)
value CERT_COMPARE_ISSUER_OF (12)
value CERT_COMPARE_KEY_IDENTIFIER (15)
value CERT_COMPARE_KEY_SPEC (9)
value CERT_COMPARE_NAME (2)
value CERT_COMPARE_NAME_STR_A (7)
value CERT_COMPARE_NAME_STR_W (8)
value CERT_COMPARE_PROPERTY (5)
value CERT_COMPARE_PUBLIC_KEY (6)
value CERT_COMPARE_SHIFT (16)
value CERT_COMPARE_SIGNATURE_HASH (14)
value CERT_COMPARE_SUBJECT_CERT (11)
value CERT_COMPARE_SUBJECT_INFO_ACCESS (19)
value CERT_CONTEXT_REVOCATION_TYPE (1)
value CERT_CREATE_SELFSIGN_NO_KEY_INFO (2)
value CERT_CREATE_SELFSIGN_NO_SIGN (1)
value CERT_CROSS_CERT_DIST_POINTS_PROP_ID (23)
value CERT_CTL_USAGE_PROP_ID (CERT_ENHKEY_USAGE_PROP_ID)
value CERT_DATE_STAMP_PROP_ID (27)
value CERT_DESCRIPTION_PROP_ID (13)
value CERT_DISALLOWED_CA_FILETIME_PROP_ID (128)
value CERT_DISALLOWED_ENHKEY_USAGE_PROP_ID (122)
value CERT_DISALLOWED_FILETIME_PROP_ID (104)
value CERT_DSS_R_LEN (20)
value CERT_DSS_S_LEN (20)
value CERT_EFS_PROP_ID (17)
value CERT_ENHKEY_USAGE_PROP_ID (9)
value CERT_ENROLLMENT_PROP_ID (26)
value CERT_EXTENDED_ERROR_INFO_PROP_ID (30)
value CERT_FILE_HASH_USE_TYPE (1)
value CERT_FIND_CTL_USAGE (CERT_FIND_ENHKEY_USAGE)
value CERT_FIND_EXT_ONLY_CTL_USAGE_FLAG (CERT_FIND_EXT_ONLY_ENHKEY_USAGE_FLAG)
value CERT_FIND_HASH (CERT_FIND_SHA1_HASH)
value CERT_FIND_ISSUER_STR (CERT_FIND_ISSUER_STR_W)
value CERT_FIND_NO_CTL_USAGE_FLAG (CERT_FIND_NO_ENHKEY_USAGE_FLAG)
value CERT_FIND_OPTIONAL_CTL_USAGE_FLAG (CERT_FIND_OPTIONAL_ENHKEY_USAGE_FLAG)
value CERT_FIND_OR_CTL_USAGE_FLAG (CERT_FIND_OR_ENHKEY_USAGE_FLAG)
value CERT_FIND_PROP_ONLY_CTL_USAGE_FLAG (CERT_FIND_PROP_ONLY_ENHKEY_USAGE_FLAG)
value CERT_FIND_SUBJECT_STR (CERT_FIND_SUBJECT_STR_W)
value CERT_FIND_VALID_CTL_USAGE_FLAG (CERT_FIND_VALID_ENHKEY_USAGE_FLAG)
value CERT_FIRST_RESERVED_PROP_ID (129)
value CERT_FORTEZZA_DATA_PROP_ID (18)
value CERT_FRIENDLY_NAME_PROP_ID (11)
value CERT_HASH_PROP_ID (CERT_SHA1_HASH_PROP_ID)
value CERT_HCRYPTPROV_OR_NCRYPT_KEY_HANDLE_PROP_ID (79)
value CERT_HCRYPTPROV_TRANSFER_PROP_ID (100)
value CERT_ID_ISSUER_SERIAL_NUMBER (1)
value CERT_ID_KEY_IDENTIFIER (2)
value CERT_INFO_EXTENSION_FLAG (11)
value CERT_INFO_ISSUER_FLAG (4)
value CERT_INFO_ISSUER_UNIQUE_ID_FLAG (9)
value CERT_INFO_NOT_AFTER_FLAG (6)
value CERT_INFO_NOT_BEFORE_FLAG (5)
value CERT_INFO_SERIAL_NUMBER_FLAG (2)
value CERT_INFO_SIGNATURE_ALGORITHM_FLAG (3)
value CERT_INFO_SUBJECT_FLAG (7)
value CERT_INFO_SUBJECT_PUBLIC_KEY_INFO_FLAG (8)
value CERT_INFO_SUBJECT_UNIQUE_ID_FLAG (10)
value CERT_INFO_VERSION_FLAG (1)
value CERT_ISOLATED_KEY_PROP_ID (118)
value CERT_ISSUER_CHAIN_PUB_KEY_CNG_ALG_BIT_LENGTH_PROP_ID (96)
value CERT_ISSUER_CHAIN_SIGN_HASH_CNG_ALG_PROP_ID (95)
value CERT_ISSUER_PUB_KEY_BIT_LENGTH_PROP_ID (94)
value CERT_KEY_CLASSIFICATION_PROP_ID (120)
value CERT_KEY_CONTEXT_PROP_ID (5)
value CERT_KEY_IDENTIFIER_PROP_ID (20)
value CERT_KEY_PROV_HANDLE_PROP_ID (1)
value CERT_KEY_PROV_INFO_PROP_ID (2)
value CERT_KEY_REPAIR_ATTEMPTED_PROP_ID (103)
value CERT_KEY_SPEC_PROP_ID (6)
value CERT_LOGOTYPE_BITS_IMAGE_RESOLUTION_CHOICE (1)
value CERT_LOGOTYPE_COLOR_IMAGE_INFO_CHOICE (2)
value CERT_LOGOTYPE_DIRECT_INFO_CHOICE (1)
value CERT_LOGOTYPE_GRAY_SCALE_IMAGE_INFO_CHOICE (1)
value CERT_LOGOTYPE_INDIRECT_INFO_CHOICE (2)
value CERT_LOGOTYPE_NO_IMAGE_RESOLUTION_CHOICE (0)
value CERT_LOGOTYPE_TABLE_SIZE_IMAGE_RESOLUTION_CHOICE (2)
value CERT_NAME_ATTR_TYPE (3)
value CERT_NAME_DNS_TYPE (6)
value CERT_NAME_EMAIL_TYPE (1)
value CERT_NAME_FRIENDLY_DISPLAY_TYPE (5)
value CERT_NAME_RDN_TYPE (2)
value CERT_NAME_SIMPLE_DISPLAY_TYPE (4)
value CERT_NAME_UPN_TYPE (8)
value CERT_NAME_URL_TYPE (7)
value CERT_NCRYPT_KEY_HANDLE_PROP_ID (78)
value CERT_NCRYPT_KEY_HANDLE_TRANSFER_PROP_ID (99)
value CERT_NEW_KEY_PROP_ID (74)
value CERT_NEXT_UPDATE_LOCATION_PROP_ID (10)
value CERT_NONCOMPLIANT_ROOT_URL_PROP_ID (123)
value CERT_NOT_BEFORE_ENHKEY_USAGE_PROP_ID (127)
value CERT_NOT_BEFORE_FILETIME_PROP_ID (126)
value CERT_NO_AUTO_EXPIRE_CHECK_PROP_ID (77)
value CERT_NO_EXPIRE_NOTIFICATION_PROP_ID (97)
value CERT_OCSP_CACHE_PREFIX_PROP_ID (75)
value CERT_OCSP_MUST_STAPLE_PROP_ID (121)
value CERT_OCSP_RESPONSE_PROP_ID (70)
value CERT_OID_NAME_STR (2)
value CERT_PUBKEY_ALG_PARA_PROP_ID (22)
value CERT_PUBKEY_HASH_RESERVED_PROP_ID (8)
value CERT_PUB_KEY_CNG_ALG_BIT_LENGTH_PROP_ID (93)
value CERT_PVK_FILE_PROP_ID (12)
value CERT_QUERY_CONTENT_CERT (1)
value CERT_QUERY_CONTENT_CERT_PAIR (13)
value CERT_QUERY_CONTENT_CRL (3)
value CERT_QUERY_CONTENT_CTL (2)
value CERT_QUERY_CONTENT_PFX (12)
value CERT_QUERY_CONTENT_PFX_AND_LOAD (14)
value CERT_QUERY_CONTENT_SERIALIZED_CERT (5)
value CERT_QUERY_CONTENT_SERIALIZED_CRL (7)
value CERT_QUERY_CONTENT_SERIALIZED_CTL (6)
value CERT_QUERY_CONTENT_SERIALIZED_STORE (4)
value CERT_QUERY_FORMAT_ASN_ASCII_HEX_ENCODED (3)
value CERT_QUERY_FORMAT_BINARY (1)
value CERT_RDN_ANY_TYPE (0)
value CERT_RDN_BMP_STRING (12)
value CERT_RDN_ENCODED_BLOB (1)
value CERT_RDN_GENERAL_STRING (10)
value CERT_RDN_GRAPHIC_STRING (8)
value CERT_RDN_NUMERIC_STRING (3)
value CERT_RDN_OCTET_STRING (2)
value CERT_RDN_PRINTABLE_STRING (4)
value CERT_RDN_TELETEX_STRING (5)
value CERT_RDN_UNICODE_STRING (12)
value CERT_RDN_UNIVERSAL_STRING (11)
value CERT_RDN_VIDEOTEX_STRING (6)
value CERT_RDN_VISIBLE_STRING (9)
value CERT_RENEWAL_PROP_ID (64)
value CERT_REQUEST_ORIGINATOR_PROP_ID (71)
value CERT_ROOT_PROGRAM_CERT_POLICIES_PROP_ID (83)
value CERT_ROOT_PROGRAM_CHAIN_POLICIES_PROP_ID (105)
value CERT_ROOT_PROGRAM_NAME_CONSTRAINTS_PROP_ID (84)
value CERT_SCARD_PIN_ID_PROP_ID (90)
value CERT_SCARD_PIN_INFO_PROP_ID (91)
value CERT_SCEP_CA_CERT_PROP_ID (111)
value CERT_SCEP_ENCRYPT_HASH_CNG_ALG_PROP_ID (114)
value CERT_SCEP_FLAGS_PROP_ID (115)
value CERT_SCEP_GUID_PROP_ID (116)
value CERT_SCEP_NONCE_PROP_ID (113)
value CERT_SCEP_RA_ENCRYPTION_CERT_PROP_ID (110)
value CERT_SCEP_RA_SIGNATURE_CERT_PROP_ID (109)
value CERT_SCEP_SERVER_CERTS_PROP_ID (108)
value CERT_SCEP_SIGNER_CERT_PROP_ID (112)
value CERT_SELECT_BY_ENHKEY_USAGE (1)
value CERT_SELECT_BY_EXTENSION (5)
value CERT_SELECT_BY_FRIENDLYNAME (13)
value CERT_SELECT_BY_ISSUER_ATTR (7)
value CERT_SELECT_BY_ISSUER_DISPLAYNAME (12)
value CERT_SELECT_BY_ISSUER_NAME (9)
value CERT_SELECT_BY_KEY_USAGE (2)
value CERT_SELECT_BY_POLICY_OID (3)
value CERT_SELECT_BY_PROV_NAME (4)
value CERT_SELECT_BY_PUBLIC_KEY (10)
value CERT_SELECT_BY_SUBJECT_ATTR (8)
value CERT_SELECT_BY_SUBJECT_HOST_NAME (6)
value CERT_SELECT_BY_THUMBPRINT (14)
value CERT_SELECT_BY_TLS_SIGNATURES (11)
value CERT_SELECT_LAST (CERT_SELECT_BY_TLS_SIGNATURES)
value CERT_SELECT_MAX_PARA (500)
value CERT_SEND_AS_TRUSTED_ISSUER_PROP_ID (102)
value CERT_SERIALIZABLE_KEY_CONTEXT_PROP_ID (117)
value CERT_SERIAL_CHAIN_PROP_ID (119)
value CERT_SIGNATURE_HASH_PROP_ID (15)
value CERT_SIGN_HASH_CNG_ALG_PROP_ID (89)
value CERT_SIMPLE_NAME_STR (1)
value CERT_SMART_CARD_DATA_PROP_ID (16)
value CERT_SMART_CARD_READER_NON_REMOVABLE_PROP_ID (106)
value CERT_SMART_CARD_READER_PROP_ID (101)
value CERT_SMART_CARD_ROOT_INFO_PROP_ID (76)
value CERT_SOURCE_LOCATION_PROP_ID (72)
value CERT_SOURCE_URL_PROP_ID (73)
value CERT_SRV_OCSP_RESP_MIN_SYNC_CERT_FILE_SECONDS_DEFAULT (5)
value CERT_STORE_ADD_ALWAYS (4)
value CERT_STORE_ADD_NEW (1)
value CERT_STORE_ADD_NEWER (6)
value CERT_STORE_ADD_NEWER_INHERIT_PROPERTIES (7)
value CERT_STORE_ADD_REPLACE_EXISTING (3)
value CERT_STORE_ADD_REPLACE_EXISTING_INHERIT_PROPERTIES (5)
value CERT_STORE_ADD_USE_EXISTING (2)
value CERT_STORE_CERTIFICATE_CONTEXT (1)
value CERT_STORE_CRL_CONTEXT (2)
value CERT_STORE_CTL_CONTEXT (3)
value CERT_STORE_CTRL_AUTO_RESYNC (4)
value CERT_STORE_CTRL_CANCEL_NOTIFY (5)
value CERT_STORE_CTRL_COMMIT (3)
value CERT_STORE_CTRL_NOTIFY_CHANGE (2)
value CERT_STORE_CTRL_RESYNC (1)
value CERT_STORE_PROV_CLOSE_FUNC (0)
value CERT_STORE_PROV_CONTROL_FUNC (13)
value CERT_STORE_PROV_DELETE_CERT_FUNC (3)
value CERT_STORE_PROV_DELETE_CRL_FUNC (7)
value CERT_STORE_PROV_DELETE_CTL_FUNC (11)
value CERT_STORE_PROV_FILENAME (CERT_STORE_PROV_FILENAME_W)
value CERT_STORE_PROV_FIND_CERT_FUNC (14)
value CERT_STORE_PROV_FIND_CRL_FUNC (17)
value CERT_STORE_PROV_FIND_CTL_FUNC (20)
value CERT_STORE_PROV_FREE_FIND_CERT_FUNC (15)
value CERT_STORE_PROV_FREE_FIND_CRL_FUNC (18)
value CERT_STORE_PROV_FREE_FIND_CTL_FUNC (21)
value CERT_STORE_PROV_GET_CERT_PROPERTY_FUNC (16)
value CERT_STORE_PROV_GET_CRL_PROPERTY_FUNC (19)
value CERT_STORE_PROV_GET_CTL_PROPERTY_FUNC (22)
value CERT_STORE_PROV_LDAP (CERT_STORE_PROV_LDAP_W)
value CERT_STORE_PROV_PHYSICAL (CERT_STORE_PROV_PHYSICAL_W)
value CERT_STORE_PROV_READ_CERT_FUNC (1)
value CERT_STORE_PROV_READ_CRL_FUNC (5)
value CERT_STORE_PROV_READ_CTL_FUNC (9)
value CERT_STORE_PROV_SET_CERT_PROPERTY_FUNC (4)
value CERT_STORE_PROV_SET_CRL_PROPERTY_FUNC (8)
value CERT_STORE_PROV_SET_CTL_PROPERTY_FUNC (12)
value CERT_STORE_PROV_SMART_CARD (CERT_STORE_PROV_SMART_CARD_W)
value CERT_STORE_PROV_SYSTEM (CERT_STORE_PROV_SYSTEM_W)
value CERT_STORE_PROV_SYSTEM_REGISTRY (CERT_STORE_PROV_SYSTEM_REGISTRY_W)
value CERT_STORE_PROV_WRITE_CERT_FUNC (2)
value CERT_STORE_PROV_WRITE_CRL_FUNC (6)
value CERT_STORE_PROV_WRITE_CTL_FUNC (10)
value CERT_STORE_SAVE_AS_STORE (1)
value CERT_STORE_SAVE_TO_FILE (1)
value CERT_STORE_SAVE_TO_FILENAME (CERT_STORE_SAVE_TO_FILENAME_W)
value CERT_STORE_SAVE_TO_FILENAME_A (3)
value CERT_STORE_SAVE_TO_FILENAME_W (4)
value CERT_STORE_SAVE_TO_MEMORY (2)
value CERT_STRONG_SIGN_OID_INFO_CHOICE (2)
value CERT_STRONG_SIGN_SERIALIZED_INFO_CHOICE (1)
value CERT_SUBJECT_DISABLE_CRL_PROP_ID (86)
value CERT_SUBJECT_INFO_ACCESS_PROP_ID (80)
value CERT_SUBJECT_OCSP_AUTHORITY_INFO_ACCESS_PROP_ID (85)
value CERT_SUBJECT_PUB_KEY_BIT_LENGTH_PROP_ID (92)
value CERT_SYSTEM_STORE_CURRENT_SERVICE_ID (4)
value CERT_SYSTEM_STORE_CURRENT_USER_GROUP_POLICY_ID (7)
value CERT_SYSTEM_STORE_CURRENT_USER_ID (1)
value CERT_SYSTEM_STORE_LOCAL_MACHINE_ENTERPRISE_ID (9)
value CERT_SYSTEM_STORE_LOCAL_MACHINE_GROUP_POLICY_ID (8)
value CERT_SYSTEM_STORE_LOCAL_MACHINE_ID (2)
value CERT_SYSTEM_STORE_LOCAL_MACHINE_WCOS_ID (10)
value CERT_SYSTEM_STORE_LOCATION_SHIFT (16)
value CERT_SYSTEM_STORE_SERVICES_ID (5)
value CERT_SYSTEM_STORE_USERS_ID (6)
value CERT_TIMESTAMP_HASH_USE_TYPE (2)
value CERT_UNICODE_ATTR_ERR_INDEX_SHIFT (16)
value CERT_UNICODE_RDN_ERR_INDEX_SHIFT (22)
value CERT_UNICODE_VALUE_ERR_INDEX_SHIFT (0)
value CERT_XML_NAME_STR (4)
value CFORCEINLINE (FORCEINLINE)
value CFSTR_MIME_NULL (NULL)
value CF_BITMAP (2)
value CF_DIB (8)
value CF_DIF (5)
value CF_ENHMETAFILE (14)
value CF_HDROP (15)
value CF_LOCALE (16)
value CF_MAX (18)
value CF_METAFILEPICT (3)
value CF_NOOEMFONTS (CF_NOVECTORFONTS)
value CF_NULL (0)
value CF_OEMTEXT (7)
value CF_PALETTE (9)
value CF_PENDATA (10)
value CF_RIFF (11)
value CF_SCRIPTSONLY (CF_ANSIONLY)
value CF_SYLK (4)
value CF_TEXT (1)
value CF_TIFF (6)
value CF_UNICODETEXT (13)
value CF_WAVE (12)
value CHAR_BIT (8)
value CHAR_MAX (SCHAR_MAX)
value CHAR_MIN (SCHAR_MIN)
value CHECKJPEGFORMAT (4119)
value CHECKPNGFORMAT (4120)
value CHILDID_SELF (0)
value CLAIM_SECURITY_ATTRIBUTES_INFORMATION_VERSION (CLAIM_SECURITY_ATTRIBUTES_INFORMATION_VERSION_V1)
value CLEARTYPE_NATURAL_QUALITY (6)
value CLEARTYPE_QUALITY (5)
value CLIPCAPS (36)
value CLIP_CHARACTER_PRECIS (1)
value CLIP_DEFAULT_PRECIS (0)
value CLIP_STROKE_PRECIS (2)
value CLIP_TO_PATH (4097)
value CLK_TCK (CLOCKS_PER_SEC)
value CLOSECHANNEL (4112)
value CLRBREAK (9)
value CLRDTR (6)
value CLRRTS (4)
value CLSID_NULL (GUID_NULL)
value CMAPI (DECLSPEC_IMPORT)
value CMC_FAIL_BAD_ALG (0)
value CMC_FAIL_BAD_CERT_ID (4)
value CMC_FAIL_BAD_IDENTITY (7)
value CMC_FAIL_BAD_MESSAGE_CHECK (1)
value CMC_FAIL_BAD_REQUEST (2)
value CMC_FAIL_BAD_TIME (3)
value CMC_FAIL_INTERNAL_CA_ERROR (11)
value CMC_FAIL_MUST_ARCHIVE_KEYS (6)
value CMC_FAIL_NO_KEY_REUSE (10)
value CMC_FAIL_POP_FAILED (9)
value CMC_FAIL_POP_REQUIRED (8)
value CMC_FAIL_TRY_LATER (12)
value CMC_FAIL_UNSUPORTED_EXT (5)
value CMC_OTHER_INFO_FAIL_CHOICE (1)
value CMC_OTHER_INFO_NO_CHOICE (0)
value CMC_OTHER_INFO_PEND_CHOICE (2)
value CMC_STATUS_CONFIRM_REQUIRED (5)
value CMC_STATUS_FAILED (2)
value CMC_STATUS_NO_SUPPORT (4)
value CMC_STATUS_PENDING (3)
value CMC_STATUS_SUCCESS (0)
value CMC_TAGGED_CERT_REQUEST_CHOICE (1)
value CMSGDATA_ALIGN (WSA_CMSGDATA_ALIGN)
value CMSGHDR_ALIGN (WSA_CMSGHDR_ALIGN)
value CMSG_ATTR_CERT_COUNT_PARAM (31)
value CMSG_ATTR_CERT_PARAM (32)
value CMSG_BARE_CONTENT_PARAM (3)
value CMSG_CERT_COUNT_PARAM (11)
value CMSG_CERT_PARAM (12)
value CMSG_CMS_RECIPIENT_COUNT_PARAM (33)
value CMSG_CMS_RECIPIENT_ENCRYPTED_KEY_INDEX_PARAM (35)
value CMSG_CMS_RECIPIENT_INDEX_PARAM (34)
value CMSG_CMS_RECIPIENT_INFO_PARAM (36)
value CMSG_CMS_SIGNER_INFO_PARAM (39)
value CMSG_COMPUTED_HASH_PARAM (22)
value CMSG_CONTENT_PARAM (2)
value CMSG_CRL_COUNT_PARAM (13)
value CMSG_CRL_PARAM (14)
value CMSG_CTRL_ADD_ATTR_CERT (14)
value CMSG_CTRL_ADD_CERT (10)
value CMSG_CTRL_ADD_CMS_SIGNER_INFO (20)
value CMSG_CTRL_ADD_CRL (12)
value CMSG_CTRL_ADD_SIGNER (6)
value CMSG_CTRL_ADD_SIGNER_UNAUTH_ATTR (8)
value CMSG_CTRL_DECRYPT (2)
value CMSG_CTRL_DEL_ATTR_CERT (15)
value CMSG_CTRL_DEL_CERT (11)
value CMSG_CTRL_DEL_CRL (13)
value CMSG_CTRL_DEL_SIGNER (7)
value CMSG_CTRL_DEL_SIGNER_UNAUTH_ATTR (9)
value CMSG_CTRL_ENABLE_STRONG_SIGNATURE (21)
value CMSG_CTRL_KEY_AGREE_DECRYPT (17)
value CMSG_CTRL_KEY_TRANS_DECRYPT (16)
value CMSG_CTRL_MAIL_LIST_DECRYPT (18)
value CMSG_CTRL_VERIFY_HASH (5)
value CMSG_CTRL_VERIFY_SIGNATURE (1)
value CMSG_CTRL_VERIFY_SIGNATURE_EX (19)
value CMSG_DATA (1)
value CMSG_ENCODED_MESSAGE (29)
value CMSG_ENCODED_SIGNER (28)
value CMSG_ENCRYPTED (6)
value CMSG_ENCRYPTED_DIGEST (27)
value CMSG_ENCRYPT_PARAM (26)
value CMSG_ENVELOPED (3)
value CMSG_ENVELOPED_DATA_CMS_VERSION (CMSG_ENVELOPED_DATA_V2)
value CMSG_ENVELOPE_ALGORITHM_PARAM (15)
value CMSG_FIRSTHDR (WSA_CMSG_FIRSTHDR)
value CMSG_HASHED (5)
value CMSG_HASHED_DATA_CMS_VERSION (CMSG_HASHED_DATA_V2)
value CMSG_HASH_ALGORITHM_PARAM (20)
value CMSG_HASH_DATA_PARAM (21)
value CMSG_INNER_CONTENT_TYPE_PARAM (4)
value CMSG_KEY_AGREE_EPHEMERAL_KEY_CHOICE (1)
value CMSG_KEY_AGREE_ORIGINATOR_CERT (1)
value CMSG_KEY_AGREE_ORIGINATOR_PUBLIC_KEY (2)
value CMSG_KEY_AGREE_RECIPIENT (2)
value CMSG_KEY_AGREE_STATIC_KEY_CHOICE (2)
value CMSG_KEY_AGREE_VERSION (CMSG_ENVELOPED_RECIPIENT_V3)
value CMSG_KEY_TRANS_CMS_VERSION (CMSG_ENVELOPED_RECIPIENT_V2)
value CMSG_KEY_TRANS_RECIPIENT (1)
value CMSG_LEN (WSA_CMSG_LEN)
value CMSG_MAIL_LIST_HANDLE_KEY_CHOICE (1)
value CMSG_MAIL_LIST_RECIPIENT (3)
value CMSG_MAIL_LIST_VERSION (CMSG_ENVELOPED_RECIPIENT_V4)
value CMSG_NXTHDR (WSA_CMSG_NXTHDR)
value CMSG_RECIPIENT_COUNT_PARAM (17)
value CMSG_RECIPIENT_INDEX_PARAM (18)
value CMSG_RECIPIENT_INFO_PARAM (19)
value CMSG_SIGNED (2)
value CMSG_SIGNED_AND_ENVELOPED (4)
value CMSG_SIGNED_DATA_CMS_VERSION (CMSG_SIGNED_DATA_V3)
value CMSG_SIGNER_AUTH_ATTR_PARAM (9)
value CMSG_SIGNER_CERT_ID_PARAM (38)
value CMSG_SIGNER_CERT_INFO_PARAM (7)
value CMSG_SIGNER_COUNT_PARAM (5)
value CMSG_SIGNER_HASH_ALGORITHM_PARAM (8)
value CMSG_SIGNER_INFO_CMS_VERSION (CMSG_SIGNER_INFO_V3)
value CMSG_SIGNER_INFO_PARAM (6)
value CMSG_SIGNER_UNAUTH_ATTR_PARAM (10)
value CMSG_SPACE (WSA_CMSG_SPACE)
value CMSG_TYPE_PARAM (1)
value CMSG_UNPROTECTED_ATTR_PARAM (37)
value CMSG_VERIFY_SIGNER_CERT (2)
value CMSG_VERIFY_SIGNER_CHAIN (3)
value CMSG_VERIFY_SIGNER_NULL (4)
value CMSG_VERIFY_SIGNER_PUBKEY (1)
value CMSG_VERSION_PARAM (30)
value CM_IN_GAMUT (0)
value CM_OUT_OF_GAMUT (255)
value CODEPAGE_ENUMPROC (CODEPAGE_ENUMPROCA)
value COLORMGMTCAPS (121)
value COLORMGMTDLGORD (1551)
value COLOROKSTRING (COLOROKSTRINGA)
value COLORONCOLOR (3)
value COLORRES (108)
value COLOR_ACTIVEBORDER (10)
value COLOR_ACTIVECAPTION (2)
value COLOR_APPWORKSPACE (12)
value COLOR_BACKGROUND (1)
value COLOR_BTNFACE (15)
value COLOR_BTNHIGHLIGHT (20)
value COLOR_BTNHILIGHT (COLOR_BTNHIGHLIGHT)
value COLOR_BTNSHADOW (16)
value COLOR_BTNTEXT (18)
value COLOR_CAPTIONTEXT (9)
value COLOR_DESKTOP (COLOR_BACKGROUND)
value COLOR_GRADIENTACTIVECAPTION (27)
value COLOR_GRADIENTINACTIVECAPTION (28)
value COLOR_GRAYTEXT (17)
value COLOR_HIGHLIGHT (13)
value COLOR_HIGHLIGHTTEXT (14)
value COLOR_HOTLIGHT (26)
value COLOR_INACTIVEBORDER (11)
value COLOR_INACTIVECAPTION (3)
value COLOR_INACTIVECAPTIONTEXT (19)
value COLOR_INFOBK (24)
value COLOR_INFOTEXT (23)
value COLOR_MENU (4)
value COLOR_MENUBAR (30)
value COLOR_MENUHILIGHT (29)
value COLOR_MENUTEXT (7)
value COLOR_SCROLLBAR (0)
value COLOR_WINDOW (5)
value COLOR_WINDOWFRAME (6)
value COLOR_WINDOWTEXT (8)
value COMPLEXREGION (3)
value COM_RIGHTS_ACTIVATE_LOCAL (8)
value COM_RIGHTS_ACTIVATE_REMOTE (16)
value COM_RIGHTS_EXECUTE (1)
value COM_RIGHTS_EXECUTE_LOCAL (2)
value COM_RIGHTS_EXECUTE_REMOTE (4)
value CONDITION_VARIABLE_INIT (RTL_CONDITION_VARIABLE_INIT)
value CONDITION_VARIABLE_LOCKMODE_SHARED (RTL_CONDITION_VARIABLE_LOCKMODE_SHARED)
value CONSOLE_FULLSCREEN (1)
value CONSOLE_FULLSCREEN_HARDWARE (2)
value CONSOLE_FULLSCREEN_MODE (1)
value CONSOLE_TEXTMODE_BUFFER (1)
value CONSOLE_WINDOWED_MODE (2)
value CONTROL_C_EXIT (STATUS_CONTROL_C_EXIT)
value CORE_PARKING_POLICY_CHANGE_IDEAL (0)
value CORE_PARKING_POLICY_CHANGE_MAX (CORE_PARKING_POLICY_CHANGE_MULTISTEP)
value CORE_PARKING_POLICY_CHANGE_MULTISTEP (3)
value CORE_PARKING_POLICY_CHANGE_ROCKET (2)
value CORE_PARKING_POLICY_CHANGE_SINGLE (1)
value CP_ACP (0)
value CP_MACCP (2)
value CP_NONE (0)
value CP_OEMCP (1)
value CP_RECTANGLE (1)
value CP_REGION (2)
value CP_SYMBOL (42)
value CP_THREAD_ACP (3)
value CP_WINANSI (1004)
value CP_WINNEUTRAL (CP_WINANSI)
value CP_WINUNICODE (1200)
value CREATE_ALWAYS (2)
value CREATE_NEW (1)
value CREATE_PROCESS_DEBUG_EVENT (3)
value CREATE_THREAD_DEBUG_EVENT (2)
value CREDENTIAL_OID_PASSWORD_CREDENTIALS (CREDENTIAL_OID_PASSWORD_CREDENTIALS_A)
value CRITICAL_SECTION_NO_DEBUG_INFO (RTL_CRITICAL_SECTION_FLAG_NO_DEBUG_INFO)
value CRL_DIST_POINT_ERR_INDEX_SHIFT (24)
value CRL_DIST_POINT_FULL_NAME (1)
value CRL_DIST_POINT_ISSUER_RDN_NAME (2)
value CRL_DIST_POINT_NO_NAME (0)
value CRL_FIND_ANY (0)
value CRL_FIND_EXISTING (2)
value CRL_FIND_ISSUED_BY (1)
value CRL_FIND_ISSUED_FOR (3)
value CRL_REASON_AA_COMPROMISE (10)
value CRL_REASON_AFFILIATION_CHANGED (3)
value CRL_REASON_CA_COMPROMISE (2)
value CRL_REASON_CERTIFICATE_HOLD (6)
value CRL_REASON_CESSATION_OF_OPERATION (5)
value CRL_REASON_KEY_COMPROMISE (1)
value CRL_REASON_PRIVILEGE_WITHDRAWN (9)
value CRL_REASON_REMOVE_FROM_CRL (8)
value CRL_REASON_SUPERSEDED (4)
value CRL_REASON_UNSPECIFIED (0)
value CROSS_CERT_DIST_POINT_ERR_INDEX_SHIFT (24)
value CRYPTNET_CACHED_OCSP_SWITCH_TO_CRL_COUNT_DEFAULT (50)
value CRYPTNET_MAX_CACHED_OCSP_PER_CRL_COUNT_DEFAULT (500)
value CRYPTNET_PRE_FETCH_AFTER_PUBLISH_PRE_FETCH_DIVISOR_DEFAULT (10)
value CRYPTNET_PRE_FETCH_BEFORE_NEXT_UPDATE_PRE_FETCH_DIVISOR_DEFAULT (20)
value CRYPTNET_PRE_FETCH_SCAN_AFTER_TRIGGER_DELAY_SECONDS_DEFAULT (60)
value CRYPTNET_PRE_FETCH_VALIDITY_PERIOD_AFTER_NEXT_UPDATE_PRE_FETCH_DIVISOR_DEFAULT (10)
value CRYPTNET_URL_CACHE_DEFAULT_FLUSH (0)
value CRYPTNET_URL_CACHE_PRE_FETCH_AUTOROOT_CAB (5)
value CRYPTNET_URL_CACHE_PRE_FETCH_BLOB (1)
value CRYPTNET_URL_CACHE_PRE_FETCH_CRL (2)
value CRYPTNET_URL_CACHE_PRE_FETCH_DISALLOWED_CERT_CAB (6)
value CRYPTNET_URL_CACHE_PRE_FETCH_NONE (0)
value CRYPTNET_URL_CACHE_PRE_FETCH_OCSP (3)
value CRYPTNET_URL_CACHE_PRE_FETCH_PIN_RULES_CAB (7)
value CRYPTNET_URL_CACHE_RESPONSE_HTTP (1)
value CRYPTNET_URL_CACHE_RESPONSE_NONE (0)
value CRYPTPROTECTMEMORY_BLOCK_SIZE (16)
value CRYPT_DEFAULT_CONTEXT_CERT_SIGN_OID (1)
value CRYPT_DEFAULT_CONTEXT_MULTI_CERT_SIGN_OID (2)
value CRYPT_DELETE_KEYSET (CRYPT_DELETEKEYSET)
value CRYPT_ECC_CMS_SHARED_INFO_SUPPPUBINFO_BYTE_LENGTH (4)
value CRYPT_ENCODE_DECODE_NONE (0)
value CRYPT_ENCRYPT_ALG_OID_GROUP_ID (2)
value CRYPT_ENHKEY_USAGE_OID_GROUP_ID (7)
value CRYPT_EXT_OR_ATTR_OID_GROUP_ID (6)
value CRYPT_FAILED (FALSE)
value CRYPT_FIRST (1)
value CRYPT_FIRST_ALG_OID_GROUP_ID (CRYPT_HASH_ALG_OID_GROUP_ID)
value CRYPT_FORMAT_CRLF (CRYPT_FORMAT_RDN_CRLF)
value CRYPT_FORMAT_SEMICOLON (CRYPT_FORMAT_RDN_SEMICOLON)
value CRYPT_HASH_ALG_OID_GROUP_ID (1)
value CRYPT_IMPL_HARDWARE (1)
value CRYPT_IMPL_MIXED (3)
value CRYPT_IMPL_REMOVABLE (8)
value CRYPT_IMPL_SOFTWARE (2)
value CRYPT_IMPL_UNKNOWN (4)
value CRYPT_INSTALL_OID_FUNC_BEFORE_FLAG (1)
value CRYPT_INSTALL_OID_INFO_BEFORE_FLAG (1)
value CRYPT_KDF_OID_GROUP_ID (10)
value CRYPT_LAST_ALG_OID_GROUP_ID (CRYPT_SIGN_ALG_OID_GROUP_ID)
value CRYPT_LAST_OID_GROUP_ID (10)
value CRYPT_LOCALIZED_NAME_ENCODING_TYPE (0)
value CRYPT_MODE_CBC (1)
value CRYPT_MODE_CBCI (6)
value CRYPT_MODE_CBCOFM (9)
value CRYPT_MODE_CBCOFMI (10)
value CRYPT_MODE_CFB (4)
value CRYPT_MODE_CFBP (7)
value CRYPT_MODE_CTS (5)
value CRYPT_MODE_ECB (2)
value CRYPT_MODE_OFB (3)
value CRYPT_MODE_OFBP (8)
value CRYPT_NEXT (2)
value CRYPT_OBJECT_LOCATOR_FIRST_RESERVED_USER_NAME_TYPE (33)
value CRYPT_OBJECT_LOCATOR_LAST_RESERVED_NAME_TYPE (32)
value CRYPT_OBJECT_LOCATOR_RELEASE_DLL_UNLOAD (4)
value CRYPT_OBJECT_LOCATOR_RELEASE_PROCESS_EXIT (3)
value CRYPT_OBJECT_LOCATOR_RELEASE_SERVICE_STOP (2)
value CRYPT_OBJECT_LOCATOR_RELEASE_SYSTEM_SHUTDOWN (1)
value CRYPT_OBJECT_LOCATOR_SPN_NAME_TYPE (1)
value CRYPT_OID_INFO_ALGID_KEY (3)
value CRYPT_OID_INFO_CNG_ALGID_KEY (5)
value CRYPT_OID_INFO_CNG_SIGN_KEY (6)
value CRYPT_OID_INFO_NAME_KEY (2)
value CRYPT_OID_INFO_OID_GROUP_BIT_LEN_SHIFT (16)
value CRYPT_OID_INFO_OID_KEY (1)
value CRYPT_OID_INFO_SIGN_KEY (4)
value CRYPT_POLICY_OID_GROUP_ID (8)
value CRYPT_PUBKEY_ALG_OID_GROUP_ID (3)
value CRYPT_RDN_ATTR_OID_GROUP_ID (5)
value CRYPT_REGISTER_FIRST_INDEX (0)
value CRYPT_SGC_ENUM (4)
value CRYPT_SIGN_ALG_OID_GROUP_ID (4)
value CRYPT_SUCCEED (TRUE)
value CRYPT_TEMPLATE_OID_GROUP_ID (9)
value CRYPT_UNICODE_NAME_ENCODE_DISABLE_CHECK_TYPE_FLAG (CERT_RDN_DISABLE_CHECK_TYPE_FLAG)
value CRYPT_USERDATA (1)
value CRYPT_VERIFY_CERT_SIGN_ISSUER_CERT (2)
value CRYPT_VERIFY_CERT_SIGN_ISSUER_CHAIN (3)
value CRYPT_VERIFY_CERT_SIGN_ISSUER_NULL (4)
value CRYPT_VERIFY_CERT_SIGN_ISSUER_PUBKEY (1)
value CRYPT_VERIFY_CERT_SIGN_SUBJECT_BLOB (1)
value CRYPT_VERIFY_CERT_SIGN_SUBJECT_CERT (2)
value CRYPT_VERIFY_CERT_SIGN_SUBJECT_CRL (3)
value CRYPT_VERIFY_CERT_SIGN_SUBJECT_OCSP_BASIC_SIGNED_RESPONSE (4)
value CSOUND_SYSTEM (16)
value CSTR_EQUAL (2)
value CSTR_GREATER_THAN (3)
value CSTR_LESS_THAN (1)
value CTLCOLOR_BTN (3)
value CTLCOLOR_DLG (4)
value CTLCOLOR_EDIT (1)
value CTLCOLOR_LISTBOX (2)
value CTLCOLOR_MAX (7)
value CTLCOLOR_MSGBOX (0)
value CTLCOLOR_SCROLLBAR (5)
value CTLCOLOR_STATIC (6)
value CTL_ANY_SUBJECT_TYPE (1)
value CTL_CERT_SUBJECT_TYPE (2)
value CTL_FIND_ANY (0)
value CTL_FIND_EXISTING (5)
value CTL_FIND_SUBJECT (4)
value CTL_FIND_USAGE (3)
value CTRL_BREAK_EVENT (1)
value CTRL_CLOSE_EVENT (2)
value CTRL_C_EVENT (0)
value CTRL_LOGOFF_EVENT (5)
value CTRL_SHUTDOWN_EVENT (6)
value CTRY_ALBANIA (355)
value CTRY_ALGERIA (213)
value CTRY_ARGENTINA (54)
value CTRY_ARMENIA (374)
value CTRY_AUSTRALIA (61)
value CTRY_AUSTRIA (43)
value CTRY_AZERBAIJAN (994)
value CTRY_BAHRAIN (973)
value CTRY_BELARUS (375)
value CTRY_BELGIUM (32)
value CTRY_BELIZE (501)
value CTRY_BOLIVIA (591)
value CTRY_BRAZIL (55)
value CTRY_BRUNEI_DARUSSALAM (673)
value CTRY_BULGARIA (359)
value CTRY_CANADA (2)
value CTRY_CARIBBEAN (1)
value CTRY_CHILE (56)
value CTRY_COLOMBIA (57)
value CTRY_COSTA_RICA (506)
value CTRY_CROATIA (385)
value CTRY_CZECH (420)
value CTRY_DEFAULT (0)
value CTRY_DENMARK (45)
value CTRY_DOMINICAN_REPUBLIC (1)
value CTRY_ECUADOR (593)
value CTRY_EGYPT (20)
value CTRY_EL_SALVADOR (503)
value CTRY_ESTONIA (372)
value CTRY_FAEROE_ISLANDS (298)
value CTRY_FINLAND (358)
value CTRY_FRANCE (33)
value CTRY_GEORGIA (995)
value CTRY_GERMANY (49)
value CTRY_GREECE (30)
value CTRY_GUATEMALA (502)
value CTRY_HONDURAS (504)
value CTRY_HONG_KONG (852)
value CTRY_HUNGARY (36)
value CTRY_ICELAND (354)
value CTRY_INDIA (91)
value CTRY_INDONESIA (62)
value CTRY_IRAN (981)
value CTRY_IRAQ (964)
value CTRY_IRELAND (353)
value CTRY_ISRAEL (972)
value CTRY_ITALY (39)
value CTRY_JAMAICA (1)
value CTRY_JAPAN (81)
value CTRY_JORDAN (962)
value CTRY_KAZAKSTAN (7)
value CTRY_KENYA (254)
value CTRY_KUWAIT (965)
value CTRY_KYRGYZSTAN (996)
value CTRY_LATVIA (371)
value CTRY_LEBANON (961)
value CTRY_LIBYA (218)
value CTRY_LIECHTENSTEIN (41)
value CTRY_LITHUANIA (370)
value CTRY_LUXEMBOURG (352)
value CTRY_MACAU (853)
value CTRY_MACEDONIA (389)
value CTRY_MALAYSIA (60)
value CTRY_MALDIVES (960)
value CTRY_MEXICO (52)
value CTRY_MONACO (33)
value CTRY_MONGOLIA (976)
value CTRY_MOROCCO (212)
value CTRY_NETHERLANDS (31)
value CTRY_NEW_ZEALAND (64)
value CTRY_NICARAGUA (505)
value CTRY_NORWAY (47)
value CTRY_OMAN (968)
value CTRY_PAKISTAN (92)
value CTRY_PANAMA (507)
value CTRY_PARAGUAY (595)
value CTRY_PERU (51)
value CTRY_PHILIPPINES (63)
value CTRY_POLAND (48)
value CTRY_PORTUGAL (351)
value CTRY_PRCHINA (86)
value CTRY_PUERTO_RICO (1)
value CTRY_QATAR (974)
value CTRY_ROMANIA (40)
value CTRY_RUSSIA (7)
value CTRY_SAUDI_ARABIA (966)
value CTRY_SERBIA (381)
value CTRY_SINGAPORE (65)
value CTRY_SLOVAK (421)
value CTRY_SLOVENIA (386)
value CTRY_SOUTH_AFRICA (27)
value CTRY_SOUTH_KOREA (82)
value CTRY_SPAIN (34)
value CTRY_SWEDEN (46)
value CTRY_SWITZERLAND (41)
value CTRY_SYRIA (963)
value CTRY_TAIWAN (886)
value CTRY_TATARSTAN (7)
value CTRY_THAILAND (66)
value CTRY_TRINIDAD_Y_TOBAGO (1)
value CTRY_TUNISIA (216)
value CTRY_TURKEY (90)
value CTRY_UAE (971)
value CTRY_UKRAINE (380)
value CTRY_UNITED_KINGDOM (44)
value CTRY_UNITED_STATES (1)
value CTRY_URUGUAY (598)
value CTRY_UZBEKISTAN (7)
value CTRY_VENEZUELA (58)
value CTRY_VIET_NAM (84)
value CTRY_YEMEN (967)
value CTRY_ZIMBABWE (263)
value CURRENT_IMPORT_REDIRECTION_VERSION (1)
value CURSOR_CREATION_SCALING_DEFAULT (2)
value CURSOR_CREATION_SCALING_NONE (1)
value CURVECAPS (28)
value CUR_BLOB_VERSION (2)
value CWCSTORAGENAME (32)
value CWMO_MAX_HANDLES (56)
value DATA_E_FORMATETC (DV_E_FORMATETC)
value DATEFMT_ENUMPROC (DATEFMT_ENUMPROCA)
value DATEFMT_ENUMPROCEX (DATEFMT_ENUMPROCEXA)
value DCB_DIRTY (DCB_ACCUMULATE)
value DCE_C_ERROR_STRING_LEN (256)
value DC_BINADJUST (19)
value DC_BINNAMES (12)
value DC_BINS (6)
value DC_BRUSH (18)
value DC_COLLATE (22)
value DC_COLORDEVICE (32)
value DC_COPIES (18)
value DC_DATATYPE_PRODUCED (21)
value DC_DRIVER (11)
value DC_DUPLEX (7)
value DC_EMF_COMPLIANT (20)
value DC_ENUMRESOLUTIONS (13)
value DC_EXTRA (9)
value DC_FIELDS (1)
value DC_FILEDEPENDENCIES (14)
value DC_MANUFACTURER (23)
value DC_MAXEXTENT (5)
value DC_MEDIAREADY (29)
value DC_MEDIATYPENAMES (34)
value DC_MEDIATYPES (35)
value DC_MINEXTENT (4)
value DC_MODEL (24)
value DC_NUP (33)
value DC_ORIENTATION (17)
value DC_PAPERNAMES (16)
value DC_PAPERS (2)
value DC_PAPERSIZE (3)
value DC_PEN (19)
value DC_PERSONALITY (25)
value DC_PRINTERMEM (28)
value DC_PRINTRATE (26)
value DC_PRINTRATEPPM (31)
value DC_PRINTRATEUNIT (27)
value DC_SIZE (8)
value DC_STAPLE (30)
value DC_TRUETYPE (15)
value DC_VERSION (10)
value DEFAULT_CHARSET (1)
value DEFAULT_GUI_FONT (17)
value DEFAULT_PALETTE (15)
value DEFAULT_PITCH (0)
value DEFAULT_QUALITY (0)
value DEF_PRIORITY (1)
value DESKTOPHORZRES (118)
value DESKTOPVERTRES (117)
value DEVICEDATA (19)
value DEVICEDUMP_MAX_IDSTRING (32)
value DEVICE_DEFAULT_FONT (14)
value DEVICE_TYPE (DWORD)
value DFC_BUTTON (4)
value DFC_CAPTION (1)
value DFC_MENU (2)
value DFC_POPUPMENU (5)
value DFC_SCROLL (3)
value DIAGNOSTIC_REASON_VERSION (0)
value DIB_PAL_COLORS (1)
value DIB_RGB_COLORS (0)
value DIFFERENCE (11)
value DISCHARGE_POLICY_CRITICAL (0)
value DISCHARGE_POLICY_LOW (1)
value DISK_BINNING (3)
value DISK_LOGGING_DUMP (2)
value DISK_LOGGING_START (0)
value DISK_LOGGING_STOP (1)
value DISPATCH_LEVEL (2)
value DISPLAYCONFIG_MAXPATH (1024)
value DISP_CHANGE_RESTART (1)
value DISP_CHANGE_SUCCESSFUL (0)
value DI_CHANNEL (1)
value DI_READ_SPOOL_JOB (3)
value DKGRAY_BRUSH (3)
value DLGWINDOWEXTRA (30)
value DLL_PROCESS_ATTACH (1)
value DLL_PROCESS_DETACH (0)
value DLL_THREAD_ATTACH (2)
value DLL_THREAD_DETACH (3)
value DMBIN_AUTO (7)
value DMBIN_CASSETTE (14)
value DMBIN_ENVELOPE (5)
value DMBIN_ENVMANUAL (6)
value DMBIN_FIRST (DMBIN_UPPER)
value DMBIN_FORMSOURCE (15)
value DMBIN_LARGECAPACITY (11)
value DMBIN_LARGEFMT (10)
value DMBIN_LAST (DMBIN_FORMSOURCE)
value DMBIN_LOWER (2)
value DMBIN_MANUAL (4)
value DMBIN_MIDDLE (3)
value DMBIN_ONLYONE (1)
value DMBIN_SMALLFMT (9)
value DMBIN_TRACTOR (8)
value DMBIN_UPPER (1)
value DMBIN_USER (256)
value DMCOLLATE_FALSE (0)
value DMCOLLATE_TRUE (1)
value DMCOLOR_COLOR (2)
value DMCOLOR_MONOCHROME (1)
value DMDFO_CENTER (2)
value DMDFO_DEFAULT (0)
value DMDFO_STRETCH (1)
value DMDITHER_COARSE (2)
value DMDITHER_ERRORDIFFUSION (5)
value DMDITHER_FINE (3)
value DMDITHER_GRAYSCALE (10)
value DMDITHER_LINEART (4)
value DMDITHER_NONE (1)
value DMDITHER_USER (256)
value DMDO_DEFAULT (0)
value DMDUP_HORIZONTAL (3)
value DMDUP_SIMPLEX (1)
value DMDUP_VERTICAL (2)
value DMICMMETHOD_DEVICE (4)
value DMICMMETHOD_DRIVER (3)
value DMICMMETHOD_NONE (1)
value DMICMMETHOD_SYSTEM (2)
value DMICMMETHOD_USER (256)
value DMICM_ABS_COLORIMETRIC (4)
value DMICM_COLORIMETRIC (3)
value DMICM_CONTRAST (2)
value DMICM_SATURATE (1)
value DMICM_USER (256)
value DMLERR_NO_ERROR (0)
value DMMEDIA_GLOSSY (3)
value DMMEDIA_STANDARD (1)
value DMMEDIA_TRANSPARENCY (2)
value DMMEDIA_USER (256)
value DMNUP_ONEUP (2)
value DMNUP_SYSTEM (1)
value DMORIENT_LANDSCAPE (2)
value DMORIENT_PORTRAIT (1)
value DMPAPER_A_PLUS (57)
value DMPAPER_B_PLUS (58)
value DMPAPER_CSHEET (24)
value DMPAPER_DBL_JAPANESE_POSTCARD (69)
value DMPAPER_DBL_JAPANESE_POSTCARD_ROTATED (82)
value DMPAPER_DSHEET (25)
value DMPAPER_ENV_DL (27)
value DMPAPER_ENV_INVITE (47)
value DMPAPER_ENV_ITALY (36)
value DMPAPER_ENV_MONARCH (37)
value DMPAPER_ENV_PERSONAL (38)
value DMPAPER_ESHEET (26)
value DMPAPER_EXECUTIVE (7)
value DMPAPER_FANFOLD_LGL_GERMAN (41)
value DMPAPER_FANFOLD_STD_GERMAN (40)
value DMPAPER_FANFOLD_US (39)
value DMPAPER_FIRST (DMPAPER_LETTER)
value DMPAPER_FOLIO (14)
value DMPAPER_JAPANESE_POSTCARD (43)
value DMPAPER_JAPANESE_POSTCARD_ROTATED (81)
value DMPAPER_LAST (DMPAPER_PENV_10_ROTATED)
value DMPAPER_LEDGER (4)
value DMPAPER_LEGAL (5)
value DMPAPER_LEGAL_EXTRA (51)
value DMPAPER_LETTER (1)
value DMPAPER_LETTERSMALL (2)
value DMPAPER_LETTER_EXTRA (50)
value DMPAPER_LETTER_EXTRA_TRANSVERSE (56)
value DMPAPER_LETTER_PLUS (59)
value DMPAPER_LETTER_ROTATED (75)
value DMPAPER_LETTER_TRANSVERSE (54)
value DMPAPER_NOTE (18)
value DMPAPER_QUARTO (15)
value DMPAPER_STATEMENT (6)
value DMPAPER_TABLOID (3)
value DMPAPER_TABLOID_EXTRA (52)
value DMPAPER_USER (256)
value DMTT_BITMAP (1)
value DMTT_DOWNLOAD (2)
value DMTT_DOWNLOAD_OUTLINE (4)
value DMTT_SUBDEV (3)
value DM_COPY (2)
value DM_IN_BUFFER (DM_MODIFY)
value DM_IN_PROMPT (DM_PROMPT)
value DM_MODIFY (8)
value DM_OUT_BUFFER (DM_COPY)
value DM_OUT_DEFAULT (DM_UPDATE)
value DM_PROMPT (4)
value DM_UPDATE (1)
value DNS_ERROR_ADDRESS_REQUIRED (9573L)
value DNS_ERROR_ALIAS_LOOP (9722L)
value DNS_ERROR_AUTOZONE_ALREADY_EXISTS (9610L)
value DNS_ERROR_AXFR (9752L)
value DNS_ERROR_BACKGROUND_LOADING (9568L)
value DNS_ERROR_BAD_KEYMASTER (9122L)
value DNS_ERROR_BAD_PACKET (9502L)
value DNS_ERROR_CANNOT_FIND_ROOT_HINTS (9564L)
value DNS_ERROR_CLIENT_SUBNET_ALREADY_EXISTS (9977L)
value DNS_ERROR_CLIENT_SUBNET_DOES_NOT_EXIST (9976L)
value DNS_ERROR_CLIENT_SUBNET_IS_ACCESSED (9975L)
value DNS_ERROR_CNAME_COLLISION (9709L)
value DNS_ERROR_CNAME_LOOP (9707L)
value DNS_ERROR_DATABASE_BASE (9700)
value DNS_ERROR_DATAFILE_BASE (9650)
value DNS_ERROR_DATAFILE_OPEN_FAILURE (9653L)
value DNS_ERROR_DATAFILE_PARSING (9655L)
value DNS_ERROR_DEFAULT_SCOPE (9960L)
value DNS_ERROR_DEFAULT_VIRTUALIZATION_INSTANCE (9925L)
value DNS_ERROR_DEFAULT_ZONESCOPE (9953L)
value DNS_ERROR_DELEGATION_REQUIRED (9571L)
value DNS_ERROR_DNAME_COLLISION (9721L)
value DNS_ERROR_DNSSEC_BASE (9100)
value DNS_ERROR_DNSSEC_IS_DISABLED (9125L)
value DNS_ERROR_DP_ALREADY_ENLISTED (9904L)
value DNS_ERROR_DP_ALREADY_EXISTS (9902L)
value DNS_ERROR_DP_BASE (9900)
value DNS_ERROR_DP_DOES_NOT_EXIST (9901L)
value DNS_ERROR_DP_FSMO_ERROR (9906L)
value DNS_ERROR_DP_NOT_AVAILABLE (9905L)
value DNS_ERROR_DP_NOT_ENLISTED (9903L)
value DNS_ERROR_DS_UNAVAILABLE (9717L)
value DNS_ERROR_DS_ZONE_ALREADY_EXISTS (9718L)
value DNS_ERROR_DWORD_VALUE_TOO_LARGE (9567L)
value DNS_ERROR_DWORD_VALUE_TOO_SMALL (9566L)
value DNS_ERROR_FILE_WRITEBACK_FAILED (9654L)
value DNS_ERROR_FORWARDER_ALREADY_EXISTS (9619L)
value DNS_ERROR_GENERAL_API_BASE (9550)
value DNS_ERROR_INCONSISTENT_ROOT_HINTS (9565L)
value DNS_ERROR_INVAILD_VIRTUALIZATION_INSTANCE_NAME (9924L)
value DNS_ERROR_INVALID_CLIENT_SUBNET_NAME (9984L)
value DNS_ERROR_INVALID_DATA (ERROR_INVALID_DATA)
value DNS_ERROR_INVALID_DATAFILE_NAME (9652L)
value DNS_ERROR_INVALID_INITIAL_ROLLOVER_OFFSET (9115L)
value DNS_ERROR_INVALID_IP_ADDRESS (9552L)
value DNS_ERROR_INVALID_KEY_SIZE (9106L)
value DNS_ERROR_INVALID_NAME (ERROR_INVALID_NAME)
value DNS_ERROR_INVALID_NAME_CHAR (9560L)
value DNS_ERROR_INVALID_POLICY_TABLE (9572L)
value DNS_ERROR_INVALID_PROPERTY (9553L)
value DNS_ERROR_INVALID_ROLLOVER_PERIOD (9114L)
value DNS_ERROR_INVALID_SCOPE_NAME (9958L)
value DNS_ERROR_INVALID_SCOPE_OPERATION (9961L)
value DNS_ERROR_INVALID_SIGNATURE_VALIDITY_PERIOD (9123L)
value DNS_ERROR_INVALID_TYPE (9551L)
value DNS_ERROR_INVALID_XML (9126L)
value DNS_ERROR_INVALID_ZONESCOPE_NAME (9954L)
value DNS_ERROR_INVALID_ZONE_OPERATION (9603L)
value DNS_ERROR_INVALID_ZONE_TYPE (9611L)
value DNS_ERROR_KEYMASTER_REQUIRED (9101L)
value DNS_ERROR_KSP_DOES_NOT_SUPPORT_PROTECTION (9108L)
value DNS_ERROR_KSP_NOT_ACCESSIBLE (9112L)
value DNS_ERROR_LOAD_ZONESCOPE_FAILED (9956L)
value DNS_ERROR_NAME_DOES_NOT_EXIST (9714L)
value DNS_ERROR_NAME_NOT_IN_ZONE (9706L)
value DNS_ERROR_NBSTAT_INIT_FAILED (9617L)
value DNS_ERROR_NEED_SECONDARY_ADDRESSES (9614L)
value DNS_ERROR_NEED_WINS_SERVERS (9616L)
value DNS_ERROR_NODE_CREATION_FAILED (9703L)
value DNS_ERROR_NODE_IS_CNAME (9708L)
value DNS_ERROR_NODE_IS_DNAME (9720L)
value DNS_ERROR_NON_RFC_NAME (9556L)
value DNS_ERROR_NOT_ALLOWED_ON_ACTIVE_SKD (9119L)
value DNS_ERROR_NOT_ALLOWED_ON_RODC (9569L)
value DNS_ERROR_NOT_ALLOWED_ON_ROOT_SERVER (9562L)
value DNS_ERROR_NOT_ALLOWED_ON_SIGNED_ZONE (9102L)
value DNS_ERROR_NOT_ALLOWED_ON_UNSIGNED_ZONE (9121L)
value DNS_ERROR_NOT_ALLOWED_ON_ZSK (9118L)
value DNS_ERROR_NOT_ALLOWED_UNDER_DELEGATION (9563L)
value DNS_ERROR_NOT_ALLOWED_UNDER_DNAME (9570L)
value DNS_ERROR_NOT_ALLOWED_WITH_ZONESCOPES (9955L)
value DNS_ERROR_NOT_ENOUGH_SIGNING_KEY_DESCRIPTORS (9104L)
value DNS_ERROR_NOT_UNIQUE (9555L)
value DNS_ERROR_NO_BOOTFILE_IF_DS_ZONE (9719L)
value DNS_ERROR_NO_CREATE_CACHE_DATA (9713L)
value DNS_ERROR_NO_DNS_SERVERS (9852L)
value DNS_ERROR_NO_MEMORY (ERROR_OUTOFMEMORY)
value DNS_ERROR_NO_PACKET (9503L)
value DNS_ERROR_NO_TCPIP (9851L)
value DNS_ERROR_NO_VALID_TRUST_ANCHORS (9127L)
value DNS_ERROR_NO_ZONE_INFO (9602L)
value DNS_ERROR_NUMERIC_NAME (9561L)
value DNS_ERROR_OPERATION_BASE (9750)
value DNS_ERROR_PACKET_FMT_BASE (9500)
value DNS_ERROR_POLICY_ALREADY_EXISTS (9971L)
value DNS_ERROR_POLICY_DOES_NOT_EXIST (9972L)
value DNS_ERROR_POLICY_INVALID_CRITERIA (9973L)
value DNS_ERROR_POLICY_INVALID_CRITERIA_CLIENT_SUBNET (9990L)
value DNS_ERROR_POLICY_INVALID_CRITERIA_FQDN (9994L)
value DNS_ERROR_POLICY_INVALID_CRITERIA_INTERFACE (9993L)
value DNS_ERROR_POLICY_INVALID_CRITERIA_NETWORK_PROTOCOL (9992L)
value DNS_ERROR_POLICY_INVALID_CRITERIA_QUERY_TYPE (9995L)
value DNS_ERROR_POLICY_INVALID_CRITERIA_TIME_OF_DAY (9996L)
value DNS_ERROR_POLICY_INVALID_CRITERIA_TRANSPORT_PROTOCOL (9991L)
value DNS_ERROR_POLICY_INVALID_NAME (9982L)
value DNS_ERROR_POLICY_INVALID_SETTINGS (9974L)
value DNS_ERROR_POLICY_INVALID_WEIGHT (9981L)
value DNS_ERROR_POLICY_LOCKED (9980L)
value DNS_ERROR_POLICY_MISSING_CRITERIA (9983L)
value DNS_ERROR_POLICY_PROCESSING_ORDER_INVALID (9985L)
value DNS_ERROR_POLICY_SCOPE_MISSING (9986L)
value DNS_ERROR_POLICY_SCOPE_NOT_ALLOWED (9987L)
value DNS_ERROR_PRIMARY_REQUIRES_DATAFILE (9651L)
value DNS_ERROR_RCODE (9504L)
value DNS_ERROR_RCODE_BADKEY (9017L)
value DNS_ERROR_RCODE_BADSIG (9016L)
value DNS_ERROR_RCODE_BADTIME (9018L)
value DNS_ERROR_RCODE_FORMAT_ERROR (9001L)
value DNS_ERROR_RCODE_LAST (DNS_ERROR_RCODE_BADTIME)
value DNS_ERROR_RCODE_NAME_ERROR (9003L)
value DNS_ERROR_RCODE_NOTAUTH (9009L)
value DNS_ERROR_RCODE_NOTZONE (9010L)
value DNS_ERROR_RCODE_NOT_IMPLEMENTED (9004L)
value DNS_ERROR_RCODE_NO_ERROR (NO_ERROR)
value DNS_ERROR_RCODE_NXRRSET (9008L)
value DNS_ERROR_RCODE_REFUSED (9005L)
value DNS_ERROR_RCODE_SERVER_FAILURE (9002L)
value DNS_ERROR_RCODE_YXDOMAIN (9006L)
value DNS_ERROR_RCODE_YXRRSET (9007L)
value DNS_ERROR_RECORD_ALREADY_EXISTS (9711L)
value DNS_ERROR_RECORD_DOES_NOT_EXIST (9701L)
value DNS_ERROR_RECORD_FORMAT (9702L)
value DNS_ERROR_RECORD_ONLY_AT_ZONE_ROOT (9710L)
value DNS_ERROR_RECORD_TIMED_OUT (9705L)
value DNS_ERROR_RESPONSE_CODES_BASE (9000)
value DNS_ERROR_ROLLOVER_ALREADY_QUEUED (9120L)
value DNS_ERROR_ROLLOVER_IN_PROGRESS (9116L)
value DNS_ERROR_ROLLOVER_NOT_POKEABLE (9128L)
value DNS_ERROR_RRL_INVALID_LEAK_RATE (9916L)
value DNS_ERROR_RRL_INVALID_TC_RATE (9915L)
value DNS_ERROR_RRL_INVALID_WINDOW_SIZE (9912L)
value DNS_ERROR_RRL_LEAK_RATE_LESSTHAN_TC_RATE (9917L)
value DNS_ERROR_RRL_NOT_ENABLED (9911L)
value DNS_ERROR_SCOPE_ALREADY_EXISTS (9963L)
value DNS_ERROR_SCOPE_DOES_NOT_EXIST (9959L)
value DNS_ERROR_SCOPE_LOCKED (9962L)
value DNS_ERROR_SECONDARY_DATA (9712L)
value DNS_ERROR_SECONDARY_REQUIRES_MASTER_IP (9612L)
value DNS_ERROR_SECURE_BASE (9800)
value DNS_ERROR_SERVERSCOPE_IS_REFERENCED (9988L)
value DNS_ERROR_SETUP_BASE (9850)
value DNS_ERROR_SIGNING_KEY_NOT_ACCESSIBLE (9107L)
value DNS_ERROR_SOA_DELETE_INVALID (9618L)
value DNS_ERROR_STANDBY_KEY_NOT_PRESENT (9117L)
value DNS_ERROR_SUBNET_ALREADY_EXISTS (9979L)
value DNS_ERROR_SUBNET_DOES_NOT_EXIST (9978L)
value DNS_ERROR_TOO_MANY_SKDS (9113L)
value DNS_ERROR_TRY_AGAIN_LATER (9554L)
value DNS_ERROR_UNEXPECTED_CNG_ERROR (9110L)
value DNS_ERROR_UNEXPECTED_DATA_PROTECTION_ERROR (9109L)
value DNS_ERROR_UNKNOWN_RECORD_TYPE (9704L)
value DNS_ERROR_UNKNOWN_SIGNING_PARAMETER_VERSION (9111L)
value DNS_ERROR_UNSECURE_PACKET (9505L)
value DNS_ERROR_UNSUPPORTED_ALGORITHM (9105L)
value DNS_ERROR_VIRTUALIZATION_INSTANCE_ALREADY_EXISTS (9921L)
value DNS_ERROR_VIRTUALIZATION_INSTANCE_DOES_NOT_EXIST (9922L)
value DNS_ERROR_VIRTUALIZATION_TREE_LOCKED (9923L)
value DNS_ERROR_WINS_INIT_FAILED (9615L)
value DNS_ERROR_ZONESCOPE_ALREADY_EXISTS (9951L)
value DNS_ERROR_ZONESCOPE_DOES_NOT_EXIST (9952L)
value DNS_ERROR_ZONESCOPE_FILE_WRITEBACK_FAILED (9957L)
value DNS_ERROR_ZONESCOPE_IS_REFERENCED (9989L)
value DNS_ERROR_ZONE_ALREADY_EXISTS (9609L)
value DNS_ERROR_ZONE_BASE (9600)
value DNS_ERROR_ZONE_CONFIGURATION_ERROR (9604L)
value DNS_ERROR_ZONE_CREATION_FAILED (9608L)
value DNS_ERROR_ZONE_DOES_NOT_EXIST (9601L)
value DNS_ERROR_ZONE_HAS_NO_NS_RECORDS (9606L)
value DNS_ERROR_ZONE_HAS_NO_SOA_RECORD (9605L)
value DNS_ERROR_ZONE_IS_SHUTDOWN (9621L)
value DNS_ERROR_ZONE_LOCKED (9607L)
value DNS_ERROR_ZONE_LOCKED_FOR_SIGNING (9622L)
value DNS_ERROR_ZONE_NOT_SECONDARY (9613L)
value DNS_ERROR_ZONE_REQUIRES_MASTER_IP (9620L)
value DNS_INFO_ADDED_LOCAL_WINS (9753L)
value DNS_INFO_AXFR_COMPLETE (9751L)
value DNS_INFO_NO_RECORDS (9501L)
value DNS_REQUEST_PENDING (9506L)
value DNS_STATUS_CONTINUE_NEEDED (9801L)
value DNS_STATUS_DOTTED_NAME (9558L)
value DNS_STATUS_FQDN (9557L)
value DNS_STATUS_PACKET_UNSECURE (DNS_ERROR_UNSECURE_PACKET)
value DNS_STATUS_SINGLE_PART_NAME (9559L)
value DNS_WARNING_DOMAIN_UNDELETED (9716L)
value DNS_WARNING_PTR_CREATE_FAILED (9715L)
value DOWNLOADFACE (514)
value DOWNLOADHEADER (4111)
value DRAFTMODE (7)
value DRAFT_QUALITY (1)
value DRAWPATTERNRECT (25)
value DRIVERVERSION (0)
value DRIVE_CDROM (5)
value DRIVE_FIXED (3)
value DRIVE_NO_ROOT_DIR (1)
value DRIVE_RAMDISK (6)
value DRIVE_REMOTE (4)
value DRIVE_REMOVABLE (2)
value DRIVE_UNKNOWN (0)
value DRV_CANCEL (DRVCNF_CANCEL)
value DRV_MCI_FIRST (DRV_RESERVED)
value DRV_OK (DRVCNF_OK)
value DRV_RESTART (DRVCNF_RESTART)
value DS_S_SUCCESS (NO_ERROR)
value DT_CHARSTREAM (4)
value DT_DISPFILE (6)
value DT_METAFILE (5)
value DT_PLOTTER (0)
value DT_RASCAMERA (3)
value DT_RASDISPLAY (1)
value DT_RASPRINTER (2)
value DWLP_MSGRESULT (0)
value EACCES (13)
value EADDRINUSE (100)
value EADDRNOTAVAIL (101)
value EAFNOSUPPORT (102)
value EAGAIN (11)
value EALREADY (103)
value EASTEUROPE_CHARSET (238)
value EBADF (9)
value EBADMSG (104)
value EBUSY (16)
value ECANCELED (105)
value ECHILD (10)
value ECONNABORTED (106)
value ECONNREFUSED (107)
value ECONNRESET (108)
value EC_DISABLE (ST_BLOCKED)
value EC_ENABLEALL (0)
value EC_ENABLEONE (ST_BLOCKNEXT)
value EC_QUERYWAITING (2)
value EDEADLK (36)
value EDEADLOCK (EDEADLK)
value EDESTADDRREQ (109)
value EDOM (33)
value EEXIST (17)
value EFAULT (14)
value EFBIG (27)
value EFS_COMPATIBILITY_VERSION_NCRYPT_PROTECTOR (5)
value EFS_COMPATIBILITY_VERSION_PFILE_PROTECTOR (6)
value EFS_EFS_SUBVER_EFS_CERT (1)
value EFS_PFILE_SUBVER_APPX (3)
value EFS_PFILE_SUBVER_RMS (2)
value EFS_SUBVER_UNKNOWN (0)
value EHOSTUNREACH (110)
value EIDRM (111)
value EILSEQ (42)
value EINPROGRESS (112)
value EINTR (4)
value EINVAL (22)
value EIO (5)
value EISCONN (113)
value EISDIR (21)
value ELF_CULTURE_LATIN (0)
value ELF_VENDOR_SIZE (4)
value ELF_VERSION (0)
value ELOOP (114)
value EMFILE (24)
value EMLINK (31)
value EMR_ABORTPATH (68)
value EMR_ALPHABLEND (114)
value EMR_ANGLEARC (41)
value EMR_ARC (45)
value EMR_ARCTO (55)
value EMR_BEGINPATH (59)
value EMR_BITBLT (76)
value EMR_CHORD (46)
value EMR_CLOSEFIGURE (61)
value EMR_COLORCORRECTPALETTE (111)
value EMR_COLORMATCHTOTARGETW (121)
value EMR_CREATEBRUSHINDIRECT (39)
value EMR_CREATECOLORSPACE (99)
value EMR_CREATECOLORSPACEW (122)
value EMR_CREATEDIBPATTERNBRUSHPT (94)
value EMR_CREATEMONOBRUSH (93)
value EMR_CREATEPALETTE (49)
value EMR_CREATEPEN (38)
value EMR_DELETECOLORSPACE (101)
value EMR_DELETEOBJECT (40)
value EMR_ELLIPSE (42)
value EMR_ENDPATH (60)
value EMR_EOF (14)
value EMR_EXCLUDECLIPRECT (29)
value EMR_EXTCREATEFONTINDIRECTW (82)
value EMR_EXTCREATEPEN (95)
value EMR_EXTFLOODFILL (53)
value EMR_EXTSELECTCLIPRGN (75)
value EMR_EXTTEXTOUTA (83)
value EMR_EXTTEXTOUTW (84)
value EMR_FILLPATH (62)
value EMR_FILLRGN (71)
value EMR_FLATTENPATH (65)
value EMR_FRAMERGN (72)
value EMR_GDICOMMENT (70)
value EMR_GLSBOUNDEDRECORD (103)
value EMR_GLSRECORD (102)
value EMR_GRADIENTFILL (118)
value EMR_HEADER (1)
value EMR_INTERSECTCLIPRECT (30)
value EMR_INVERTRGN (73)
value EMR_LINETO (54)
value EMR_MASKBLT (78)
value EMR_MAX (122)
value EMR_MIN (1)
value EMR_MODIFYWORLDTRANSFORM (36)
value EMR_MOVETOEX (27)
value EMR_OFFSETCLIPRGN (26)
value EMR_PAINTRGN (74)
value EMR_PIE (47)
value EMR_PIXELFORMAT (104)
value EMR_PLGBLT (79)
value EMR_POLYBEZIER (2)
value EMR_POLYBEZIERTO (5)
value EMR_POLYDRAW (56)
value EMR_POLYGON (3)
value EMR_POLYLINE (4)
value EMR_POLYLINETO (6)
value EMR_POLYPOLYGON (8)
value EMR_POLYPOLYLINE (7)
value EMR_POLYTEXTOUTA (96)
value EMR_POLYTEXTOUTW (97)
value EMR_REALIZEPALETTE (52)
value EMR_RECTANGLE (43)
value EMR_RESIZEPALETTE (51)
value EMR_RESTOREDC (34)
value EMR_ROUNDRECT (44)
value EMR_SAVEDC (33)
value EMR_SCALEVIEWPORTEXTEX (31)
value EMR_SCALEWINDOWEXTEX (32)
value EMR_SELECTCLIPPATH (67)
value EMR_SELECTOBJECT (37)
value EMR_SELECTPALETTE (48)
value EMR_SETARCDIRECTION (57)
value EMR_SETBKCOLOR (25)
value EMR_SETBKMODE (18)
value EMR_SETBRUSHORGEX (13)
value EMR_SETCOLORADJUSTMENT (23)
value EMR_SETCOLORSPACE (100)
value EMR_SETDIBITSTODEVICE (80)
value EMR_SETICMMODE (98)
value EMR_SETICMPROFILEA (112)
value EMR_SETICMPROFILEW (113)
value EMR_SETLAYOUT (115)
value EMR_SETMAPMODE (17)
value EMR_SETMAPPERFLAGS (16)
value EMR_SETMETARGN (28)
value EMR_SETMITERLIMIT (58)
value EMR_SETPALETTEENTRIES (50)
value EMR_SETPIXELV (15)
value EMR_SETPOLYFILLMODE (19)
value EMR_SETSTRETCHBLTMODE (21)
value EMR_SETTEXTALIGN (22)
value EMR_SETTEXTCOLOR (24)
value EMR_SETVIEWPORTEXTEX (11)
value EMR_SETVIEWPORTORGEX (12)
value EMR_SETWINDOWEXTEX (9)
value EMR_SETWINDOWORGEX (10)
value EMR_SETWORLDTRANSFORM (35)
value EMR_STRETCHBLT (77)
value EMR_STRETCHDIBITS (81)
value EMR_STROKEANDFILLPATH (63)
value EMR_STROKEPATH (64)
value EMR_TRANSPARENTBLT (116)
value EMR_WIDENPATH (66)
value EMSGSIZE (115)
value EM_SETLIMITTEXT (EM_LIMITTEXT)
value ENABLEDUPLEX (28)
value ENABLEPAIRKERNING (769)
value ENABLERELATIVEWIDTHS (768)
value ENAMETOOLONG (38)
value ENCAPSULATED_POSTSCRIPT (4116)
value ENCLAVE_LONG_ID_LENGTH (32)
value ENCLAVE_SHORT_ID_LENGTH (16)
value ENCRYPTED_DATA_INFO_SPARSE_FILE (1)
value ENDDOC (11)
value END_PATH (4098)
value ENETDOWN (116)
value ENETRESET (117)
value ENETUNREACH (118)
value ENFILE (23)
value ENOBUFS (119)
value ENODATA (120)
value ENODEV (19)
value ENOENT (2)
value ENOEXEC (8)
value ENOLCK (39)
value ENOLINK (121)
value ENOMEM (12)
value ENOMSG (122)
value ENOPROTOOPT (123)
value ENOSPC (28)
value ENOSR (124)
value ENOSTR (125)
value ENOSYS (40)
value ENOTCONN (126)
value ENOTDIR (20)
value ENOTEMPTY (41)
value ENOTRECOVERABLE (127)
value ENOTSOCK (128)
value ENOTSUP (129)
value ENOTTY (25)
value ENUMPAPERBINS (31)
value ENUMPAPERMETRICS (34)
value ENUMRESLANGPROC (ENUMRESLANGPROCA)
value ENUMRESNAMEPROC (ENUMRESNAMEPROCA)
value ENUMRESTYPEPROC (ENUMRESTYPEPROCA)
value ENXIO (6)
value EOPNOTSUPP (130)
value EOTHER (131)
value EOVERFLOW (132)
value EOWNERDEAD (133)
value EPERM (1)
value EPIPE (32)
value EPROTO (134)
value EPROTONOSUPPORT (135)
value EPROTOTYPE (136)
value EPSPRINTING (33)
value EPT_S_CANT_CREATE (1899L)
value EPT_S_CANT_PERFORM_OP (1752L)
value EPT_S_INVALID_ENTRY (1751L)
value EPT_S_NOT_REGISTERED (1753L)
value ERANGE (34)
value EROFS (30)
value ERROR (0)
value ERROR_ABANDON_HIBERFILE (787L)
value ERROR_ABIOS_ERROR (538L)
value ERROR_ACCESS_AUDIT_BY_POLICY (785L)
value ERROR_ACCESS_DENIED (5L)
value ERROR_ACCESS_DENIED_APPDATA (502L)
value ERROR_ACCESS_DISABLED_BY_POLICY (1260L)
value ERROR_ACCESS_DISABLED_NO_SAFER_UI_BY_POLICY (786L)
value ERROR_ACCESS_DISABLED_WEBBLADE (1277L)
value ERROR_ACCESS_DISABLED_WEBBLADE_TAMPER (1278L)
value ERROR_ACCOUNT_DISABLED (1331L)
value ERROR_ACCOUNT_EXPIRED (1793L)
value ERROR_ACCOUNT_LOCKED_OUT (1909L)
value ERROR_ACCOUNT_RESTRICTION (1327L)
value ERROR_ACPI_ERROR (669L)
value ERROR_ACTIVATION_COUNT_EXCEEDED (7059L)
value ERROR_ACTIVE_CONNECTIONS (2402L)
value ERROR_ADAP_HDW_ERR (57L)
value ERROR_ADDRESS_ALREADY_ASSOCIATED (1227L)
value ERROR_ADDRESS_NOT_ASSOCIATED (1228L)
value ERROR_ADVANCED_INSTALLER_FAILED (14099L)
value ERROR_ALERTED (739L)
value ERROR_ALIAS_EXISTS (1379L)
value ERROR_ALLOCATE_BUCKET (602L)
value ERROR_ALLOTTED_SPACE_EXCEEDED (1344L)
value ERROR_ALL_NODES_NOT_AVAILABLE (5037L)
value ERROR_ALL_USER_TRUST_QUOTA_EXCEEDED (1933L)
value ERROR_ALREADY_ASSIGNED (85L)
value ERROR_ALREADY_EXISTS (183L)
value ERROR_ALREADY_FIBER (1280L)
value ERROR_ALREADY_HAS_STREAM_ID (4444L)
value ERROR_ALREADY_INITIALIZED (1247L)
value ERROR_ALREADY_REGISTERED (1242L)
value ERROR_ALREADY_RUNNING_LKG (1074L)
value ERROR_ALREADY_THREAD (1281L)
value ERROR_ALREADY_WAITING (1904L)
value ERROR_AMBIGUOUS_SYSTEM_DEVICE (15250L)
value ERROR_API_UNAVAILABLE (15841L)
value ERROR_APPCONTAINER_REQUIRED (4251L)
value ERROR_APPEXEC_APP_COMPAT_BLOCK (3068L)
value ERROR_APPEXEC_CALLER_WAIT_TIMEOUT (3069L)
value ERROR_APPEXEC_CALLER_WAIT_TIMEOUT_LICENSING (3071L)
value ERROR_APPEXEC_CALLER_WAIT_TIMEOUT_RESOURCES (3072L)
value ERROR_APPEXEC_CALLER_WAIT_TIMEOUT_TERMINATION (3070L)
value ERROR_APPEXEC_CONDITION_NOT_SATISFIED (3060L)
value ERROR_APPEXEC_HANDLE_INVALIDATED (3061L)
value ERROR_APPEXEC_HOST_ID_MISMATCH (3066L)
value ERROR_APPEXEC_INVALID_HOST_GENERATION (3062L)
value ERROR_APPEXEC_INVALID_HOST_STATE (3064L)
value ERROR_APPEXEC_NO_DONOR (3065L)
value ERROR_APPEXEC_UNEXPECTED_PROCESS_REGISTRATION (3063L)
value ERROR_APPEXEC_UNKNOWN_USER (3067L)
value ERROR_APPHELP_BLOCK (1259L)
value ERROR_APPINSTALLER_ACTIVATION_BLOCKED (15646L)
value ERROR_APPINSTALLER_IS_MANAGED_BY_SYSTEM (15672L)
value ERROR_APPINSTALLER_URI_IN_USE (15671L)
value ERROR_APPX_FILE_NOT_ENCRYPTED (409L)
value ERROR_APPX_INTEGRITY_FAILURE_CLR_NGEN (15624L)
value ERROR_APPX_RAW_DATA_WRITE_FAILED (15648L)
value ERROR_APP_DATA_CORRUPT (4402L)
value ERROR_APP_DATA_EXPIRED (4401L)
value ERROR_APP_DATA_LIMIT_EXCEEDED (4403L)
value ERROR_APP_DATA_NOT_FOUND (4400L)
value ERROR_APP_DATA_REBOOT_REQUIRED (4404L)
value ERROR_APP_HANG (1298L)
value ERROR_APP_INIT_FAILURE (575L)
value ERROR_APP_WRONG_OS (1151L)
value ERROR_ARBITRATION_UNHANDLED (723L)
value ERROR_ARENA_TRASHED (7L)
value ERROR_ARITHMETIC_OVERFLOW (534L)
value ERROR_ASSERTION_FAILURE (668L)
value ERROR_ATOMIC_LOCKS_NOT_SUPPORTED (174L)
value ERROR_AUDIT_FAILED (606L)
value ERROR_AUTHENTICATION_FIREWALL_FAILED (1935L)
value ERROR_AUTHIP_FAILURE (1469L)
value ERROR_BACKUP_CONTROLLER (586L)
value ERROR_BADDB (1009L)
value ERROR_BADKEY (1010L)
value ERROR_BADSTARTPOSITION (778L)
value ERROR_BAD_ACCESSOR_FLAGS (773L)
value ERROR_BAD_ARGUMENTS (160L)
value ERROR_BAD_CLUSTERS (6849L)
value ERROR_BAD_COMMAND (22L)
value ERROR_BAD_COMPRESSION_BUFFER (605L)
value ERROR_BAD_CONFIGURATION (1610L)
value ERROR_BAD_CURRENT_DIRECTORY (703L)
value ERROR_BAD_DESCRIPTOR_FORMAT (1361L)
value ERROR_BAD_DEVICE (1200L)
value ERROR_BAD_DEVICE_PATH (330L)
value ERROR_BAD_DEV_TYPE (66L)
value ERROR_BAD_DLL_ENTRYPOINT (609L)
value ERROR_BAD_DRIVER (2001L)
value ERROR_BAD_DRIVER_LEVEL (119L)
value ERROR_BAD_ENVIRONMENT (10L)
value ERROR_BAD_EXE_FORMAT (193L)
value ERROR_BAD_FILE_TYPE (222L)
value ERROR_BAD_FORMAT (11L)
value ERROR_BAD_FUNCTION_TABLE (559L)
value ERROR_BAD_IMPERSONATION_LEVEL (1346L)
value ERROR_BAD_INHERITANCE_ACL (1340L)
value ERROR_BAD_LENGTH (24L)
value ERROR_BAD_LOGON_SESSION_STATE (1365L)
value ERROR_BAD_MCFG_TABLE (791L)
value ERROR_BAD_NETPATH (53L)
value ERROR_BAD_NET_NAME (67L)
value ERROR_BAD_NET_RESP (58L)
value ERROR_BAD_PATHNAME (161L)
value ERROR_BAD_PIPE (230L)
value ERROR_BAD_PROFILE (1206L)
value ERROR_BAD_PROVIDER (1204L)
value ERROR_BAD_QUERY_SYNTAX (1615L)
value ERROR_BAD_RECOVERY_POLICY (6012L)
value ERROR_BAD_REM_ADAP (60L)
value ERROR_BAD_SERVICE_ENTRYPOINT (610L)
value ERROR_BAD_STACK (543L)
value ERROR_BAD_THREADID_ADDR (159L)
value ERROR_BAD_TOKEN_TYPE (1349L)
value ERROR_BAD_UNIT (20L)
value ERROR_BAD_USERNAME (2202L)
value ERROR_BAD_USER_PROFILE (1253L)
value ERROR_BAD_VALIDATION_CLASS (1348L)
value ERROR_BEGINNING_OF_MEDIA (1102L)
value ERROR_BEYOND_VDL (1289L)
value ERROR_BIDI_ERROR_BASE (13000)
value ERROR_BIDI_NOT_SUPPORTED (ERROR_NOT_SUPPORTED)
value ERROR_BIDI_STATUS_OK (0)
value ERROR_BIOS_FAILED_TO_CONNECT_INTERRUPT (585L)
value ERROR_BLOCKED_BY_PARENTAL_CONTROLS (346L)
value ERROR_BLOCK_SHARED (514L)
value ERROR_BLOCK_SOURCE_WEAK_REFERENCE_INVALID (512L)
value ERROR_BLOCK_TARGET_WEAK_REFERENCE_INVALID (513L)
value ERROR_BLOCK_TOO_MANY_REFERENCES (347L)
value ERROR_BLOCK_WEAK_REFERENCE_INVALID (511L)
value ERROR_BOOT_ALREADY_ACCEPTED (1076L)
value ERROR_BROKEN_PIPE (109L)
value ERROR_BUFFER_ALL_ZEROS (754L)
value ERROR_BUFFER_OVERFLOW (111L)
value ERROR_BUSY (170L)
value ERROR_BUSY_DRIVE (142L)
value ERROR_BUS_RESET (1111L)
value ERROR_BYPASSIO_FLT_NOT_SUPPORTED (506L)
value ERROR_CACHE_PAGE_LOCKED (752L)
value ERROR_CALLBACK_INVOKE_INLINE (812L)
value ERROR_CALLBACK_POP_STACK (768L)
value ERROR_CALLBACK_SUPPLIED_INVALID_DATA (1273L)
value ERROR_CALL_NOT_IMPLEMENTED (120L)
value ERROR_CANCELLED (1223L)
value ERROR_CANCEL_VIOLATION (173L)
value ERROR_CANNOT_ABORT_TRANSACTIONS (6848L)
value ERROR_CANNOT_ACCEPT_TRANSACTED_WORK (6847L)
value ERROR_CANNOT_BREAK_OPLOCK (802L)
value ERROR_CANNOT_COPY (266L)
value ERROR_CANNOT_DETECT_DRIVER_FAILURE (1080L)
value ERROR_CANNOT_DETECT_PROCESS_ABORT (1081L)
value ERROR_CANNOT_EXECUTE_FILE_IN_TRANSACTION (6838L)
value ERROR_CANNOT_FIND_WND_CLASS (1407L)
value ERROR_CANNOT_GRANT_REQUESTED_OPLOCK (801L)
value ERROR_CANNOT_IMPERSONATE (1368L)
value ERROR_CANNOT_LOAD_REGISTRY_FILE (589L)
value ERROR_CANNOT_MAKE (82L)
value ERROR_CANNOT_OPEN_PROFILE (1205L)
value ERROR_CANNOT_SWITCH_RUNLEVEL (15400L)
value ERROR_CANTFETCHBACKWARDS (770L)
value ERROR_CANTOPEN (1011L)
value ERROR_CANTREAD (1012L)
value ERROR_CANTSCROLLBACKWARDS (771L)
value ERROR_CANTWRITE (1013L)
value ERROR_CANT_ACCESS_DOMAIN_INFO (1351L)
value ERROR_CANT_ACCESS_FILE (1920L)
value ERROR_CANT_BREAK_TRANSACTIONAL_DEPENDENCY (6824L)
value ERROR_CANT_CLEAR_ENCRYPTION_FLAG (432L)
value ERROR_CANT_CREATE_MORE_STREAM_MINIVERSIONS (6812L)
value ERROR_CANT_CROSS_RM_BOUNDARY (6825L)
value ERROR_CANT_DELETE_LAST_ITEM (4335L)
value ERROR_CANT_DISABLE_MANDATORY (1310L)
value ERROR_CANT_ENABLE_DENY_ONLY (629L)
value ERROR_CANT_EVICT_ACTIVE_NODE (5009L)
value ERROR_CANT_OPEN_ANONYMOUS (1347L)
value ERROR_CANT_OPEN_MINIVERSION_WITH_MODIFY_INTENT (6811L)
value ERROR_CANT_RECOVER_WITH_HANDLE_OPEN (6818L)
value ERROR_CANT_RESOLVE_FILENAME (1921L)
value ERROR_CANT_TERMINATE_SELF (555L)
value ERROR_CANT_WAIT (554L)
value ERROR_CAN_NOT_COMPLETE (1003L)
value ERROR_CAN_NOT_DEL_LOCAL_WINS (4001L)
value ERROR_CAPAUTHZ_CHANGE_TYPE (451L)
value ERROR_CAPAUTHZ_DB_CORRUPTED (455L)
value ERROR_CAPAUTHZ_NOT_AUTHORIZED (453L)
value ERROR_CAPAUTHZ_NOT_DEVUNLOCKED (450L)
value ERROR_CAPAUTHZ_NOT_PROVISIONED (452L)
value ERROR_CAPAUTHZ_NO_POLICY (454L)
value ERROR_CAPAUTHZ_SCCD_DEV_MODE_REQUIRED (459L)
value ERROR_CAPAUTHZ_SCCD_INVALID_CATALOG (456L)
value ERROR_CAPAUTHZ_SCCD_NO_AUTH_ENTITY (457L)
value ERROR_CAPAUTHZ_SCCD_NO_CAPABILITY_MATCH (460L)
value ERROR_CAPAUTHZ_SCCD_PARSE_ERROR (458L)
value ERROR_CARDBUS_NOT_SUPPORTED (724L)
value ERROR_CASE_DIFFERING_NAMES_IN_DIR (424L)
value ERROR_CASE_SENSITIVE_PATH (442L)
value ERROR_CERTIFICATE_VALIDATION_PREFERENCE_CONFLICT (817L)
value ERROR_CHECKING_FILE_SYSTEM (712L)
value ERROR_CHECKOUT_REQUIRED (221L)
value ERROR_CHILD_MUST_BE_VOLATILE (1021L)
value ERROR_CHILD_NOT_COMPLETE (129L)
value ERROR_CHILD_PROCESS_BLOCKED (367L)
value ERROR_CHILD_WINDOW_MENU (1436L)
value ERROR_CIMFS_IMAGE_CORRUPT (470L)
value ERROR_CIMFS_IMAGE_VERSION_NOT_SUPPORTED (471L)
value ERROR_CIRCULAR_DEPENDENCY (1059L)
value ERROR_CLASSIC_COMPAT_MODE_NOT_ALLOWED (15667L)
value ERROR_CLASS_ALREADY_EXISTS (1410L)
value ERROR_CLASS_DOES_NOT_EXIST (1411L)
value ERROR_CLASS_HAS_WINDOWS (1412L)
value ERROR_CLEANER_CARTRIDGE_INSTALLED (4340L)
value ERROR_CLEANER_CARTRIDGE_SPENT (4333L)
value ERROR_CLEANER_SLOT_NOT_SET (4332L)
value ERROR_CLEANER_SLOT_SET (4331L)
value ERROR_CLIENT_SERVER_PARAMETERS_INVALID (597L)
value ERROR_CLIPBOARD_NOT_OPEN (1418L)
value ERROR_CLIPPING_NOT_SUPPORTED (2005L)
value ERROR_CLOUD_FILE_ACCESS_DENIED (395L)
value ERROR_CLOUD_FILE_ALREADY_CONNECTED (378L)
value ERROR_CLOUD_FILE_AUTHENTICATION_FAILED (386L)
value ERROR_CLOUD_FILE_CONNECTED_PROVIDER_ONLY (382L)
value ERROR_CLOUD_FILE_DEHYDRATION_DISALLOWED (434L)
value ERROR_CLOUD_FILE_INCOMPATIBLE_HARDLINKS (396L)
value ERROR_CLOUD_FILE_INSUFFICIENT_RESOURCES (387L)
value ERROR_CLOUD_FILE_INVALID_REQUEST (380L)
value ERROR_CLOUD_FILE_IN_USE (391L)
value ERROR_CLOUD_FILE_METADATA_CORRUPT (363L)
value ERROR_CLOUD_FILE_METADATA_TOO_LARGE (364L)
value ERROR_CLOUD_FILE_NETWORK_UNAVAILABLE (388L)
value ERROR_CLOUD_FILE_NOT_IN_SYNC (377L)
value ERROR_CLOUD_FILE_NOT_SUPPORTED (379L)
value ERROR_CLOUD_FILE_NOT_UNDER_SYNC_ROOT (390L)
value ERROR_CLOUD_FILE_PINNED (392L)
value ERROR_CLOUD_FILE_PROPERTY_BLOB_CHECKSUM_MISMATCH (366L)
value ERROR_CLOUD_FILE_PROPERTY_BLOB_TOO_LARGE (365L)
value ERROR_CLOUD_FILE_PROPERTY_CORRUPT (394L)
value ERROR_CLOUD_FILE_PROPERTY_LOCK_CONFLICT (397L)
value ERROR_CLOUD_FILE_PROPERTY_VERSION_NOT_SUPPORTED (375L)
value ERROR_CLOUD_FILE_PROVIDER_NOT_RUNNING (362L)
value ERROR_CLOUD_FILE_PROVIDER_TERMINATED (404L)
value ERROR_CLOUD_FILE_READ_ONLY_VOLUME (381L)
value ERROR_CLOUD_FILE_REQUEST_ABORTED (393L)
value ERROR_CLOUD_FILE_REQUEST_CANCELED (398L)
value ERROR_CLOUD_FILE_REQUEST_TIMEOUT (426L)
value ERROR_CLOUD_FILE_SYNC_ROOT_METADATA_CORRUPT (358L)
value ERROR_CLOUD_FILE_TOO_MANY_PROPERTY_BLOBS (374L)
value ERROR_CLOUD_FILE_UNSUCCESSFUL (389L)
value ERROR_CLOUD_FILE_US_MESSAGE_TIMEOUT (475L)
value ERROR_CLOUD_FILE_VALIDATION_FAILED (383L)
value ERROR_CLUSCFG_ALREADY_COMMITTED (5901L)
value ERROR_CLUSCFG_ROLLBACK_FAILED (5902L)
value ERROR_CLUSCFG_SYSTEM_DISK_DRIVE_LETTER_CONFLICT (5903L)
value ERROR_CLUSTERLOG_CHKPOINT_NOT_FOUND (5032L)
value ERROR_CLUSTERLOG_CORRUPT (5029L)
value ERROR_CLUSTERLOG_EXCEEDS_MAXSIZE (5031L)
value ERROR_CLUSTERLOG_NOT_ENOUGH_SPACE (5033L)
value ERROR_CLUSTERLOG_RECORD_EXCEEDS_MAXSIZE (5030L)
value ERROR_CLUSTERSET_MANAGEMENT_CLUSTER_UNREACHABLE (5999L)
value ERROR_CLUSTER_AFFINITY_CONFLICT (5971L)
value ERROR_CLUSTER_BACKUP_IN_PROGRESS (5949L)
value ERROR_CLUSTER_CANNOT_RETURN_PROPERTIES (5968L)
value ERROR_CLUSTER_CANT_CREATE_DUP_CLUSTER_NAME (5900L)
value ERROR_CLUSTER_CANT_DESERIALIZE_DATA (5923L)
value ERROR_CLUSTER_CSV_INVALID_HANDLE (5989L)
value ERROR_CLUSTER_CSV_IO_PAUSE_TIMEOUT (5979L)
value ERROR_CLUSTER_CSV_SUPPORTED_ONLY_ON_COORDINATOR (5990L)
value ERROR_CLUSTER_DATABASE_SEQMISMATCH (5083L)
value ERROR_CLUSTER_DATABASE_TRANSACTION_IN_PROGRESS (5918L)
value ERROR_CLUSTER_DATABASE_TRANSACTION_NOT_IN_PROGRESS (5919L)
value ERROR_CLUSTER_DATABASE_UPDATE_CONDITION_FAILED (5986L)
value ERROR_CLUSTER_DISK_NOT_CONNECTED (5963L)
value ERROR_CLUSTER_EVICT_INVALID_REQUEST (5939L)
value ERROR_CLUSTER_EVICT_WITHOUT_CLEANUP (5896L)
value ERROR_CLUSTER_FAULT_DOMAIN_INVALID_HIERARCHY (5995L)
value ERROR_CLUSTER_FAULT_DOMAIN_PARENT_NOT_FOUND (5994L)
value ERROR_CLUSTER_GROUP_BUSY (5944L)
value ERROR_CLUSTER_GROUP_MOVING (5908L)
value ERROR_CLUSTER_GROUP_QUEUED (5959L)
value ERROR_CLUSTER_GROUP_SINGLETON_RESOURCE (5941L)
value ERROR_CLUSTER_GUM_NOT_LOCKER (5085L)
value ERROR_CLUSTER_INCOMPATIBLE_VERSIONS (5075L)
value ERROR_CLUSTER_INSTANCE_ID_MISMATCH (5893L)
value ERROR_CLUSTER_INTERNAL_INVALID_FUNCTION (5912L)
value ERROR_CLUSTER_INVALID_INFRASTRUCTURE_FILESERVER_NAME (5998L)
value ERROR_CLUSTER_INVALID_NETWORK (5054L)
value ERROR_CLUSTER_INVALID_NETWORK_PROVIDER (5049L)
value ERROR_CLUSTER_INVALID_NODE (5039L)
value ERROR_CLUSTER_INVALID_NODE_WEIGHT (5954L)
value ERROR_CLUSTER_INVALID_REQUEST (5048L)
value ERROR_CLUSTER_INVALID_SECURITY_DESCRIPTOR (5946L)
value ERROR_CLUSTER_INVALID_STRING_FORMAT (5917L)
value ERROR_CLUSTER_INVALID_STRING_TERMINATION (5916L)
value ERROR_CLUSTER_IPADDR_IN_USE (5057L)
value ERROR_CLUSTER_JOIN_ABORTED (5074L)
value ERROR_CLUSTER_JOIN_IN_PROGRESS (5041L)
value ERROR_CLUSTER_JOIN_NOT_IN_PROGRESS (5053L)
value ERROR_CLUSTER_LAST_INTERNAL_NETWORK (5066L)
value ERROR_CLUSTER_LOCAL_NODE_NOT_FOUND (5043L)
value ERROR_CLUSTER_MAXNUM_OF_RESOURCES_EXCEEDED (5076L)
value ERROR_CLUSTER_MAX_NODES_IN_CLUSTER (5934L)
value ERROR_CLUSTER_MEMBERSHIP_HALT (5892L)
value ERROR_CLUSTER_MEMBERSHIP_INVALID_STATE (5890L)
value ERROR_CLUSTER_MISMATCHED_COMPUTER_ACCT_NAME (5905L)
value ERROR_CLUSTER_NETINTERFACE_EXISTS (5046L)
value ERROR_CLUSTER_NETINTERFACE_NOT_FOUND (5047L)
value ERROR_CLUSTER_NETWORK_ALREADY_OFFLINE (5064L)
value ERROR_CLUSTER_NETWORK_ALREADY_ONLINE (5063L)
value ERROR_CLUSTER_NETWORK_EXISTS (5044L)
value ERROR_CLUSTER_NETWORK_HAS_DEPENDENTS (5067L)
value ERROR_CLUSTER_NETWORK_NOT_FOUND (5045L)
value ERROR_CLUSTER_NETWORK_NOT_FOUND_FOR_IP (5894L)
value ERROR_CLUSTER_NETWORK_NOT_INTERNAL (5060L)
value ERROR_CLUSTER_NODE_ALREADY_DOWN (5062L)
value ERROR_CLUSTER_NODE_ALREADY_HAS_DFS_ROOT (5088L)
value ERROR_CLUSTER_NODE_ALREADY_MEMBER (5065L)
value ERROR_CLUSTER_NODE_ALREADY_UP (5061L)
value ERROR_CLUSTER_NODE_DOWN (5050L)
value ERROR_CLUSTER_NODE_DRAIN_IN_PROGRESS (5962L)
value ERROR_CLUSTER_NODE_EXISTS (5040L)
value ERROR_CLUSTER_NODE_IN_GRACE_PERIOD (5978L)
value ERROR_CLUSTER_NODE_ISOLATED (5984L)
value ERROR_CLUSTER_NODE_NOT_FOUND (5042L)
value ERROR_CLUSTER_NODE_NOT_MEMBER (5052L)
value ERROR_CLUSTER_NODE_NOT_PAUSED (5058L)
value ERROR_CLUSTER_NODE_NOT_READY (5072L)
value ERROR_CLUSTER_NODE_PAUSED (5070L)
value ERROR_CLUSTER_NODE_QUARANTINED (5985L)
value ERROR_CLUSTER_NODE_SHUTTING_DOWN (5073L)
value ERROR_CLUSTER_NODE_UNREACHABLE (5051L)
value ERROR_CLUSTER_NODE_UP (5056L)
value ERROR_CLUSTER_NOT_INSTALLED (5932L)
value ERROR_CLUSTER_NOT_SHARED_VOLUME (5945L)
value ERROR_CLUSTER_NO_NET_ADAPTERS (5906L)
value ERROR_CLUSTER_NO_QUORUM (5925L)
value ERROR_CLUSTER_NO_RPC_PACKAGES_REGISTERED (5081L)
value ERROR_CLUSTER_NO_SECURITY_CONTEXT (5059L)
value ERROR_CLUSTER_NULL_DATA (5920L)
value ERROR_CLUSTER_OBJECT_ALREADY_USED (5936L)
value ERROR_CLUSTER_OBJECT_IS_CLUSTER_SET_VM (6250L)
value ERROR_CLUSTER_OLD_VERSION (5904L)
value ERROR_CLUSTER_OWNER_NOT_IN_PREFLIST (5082L)
value ERROR_CLUSTER_PARAMETER_MISMATCH (5897L)
value ERROR_CLUSTER_PARAMETER_OUT_OF_BOUNDS (5913L)
value ERROR_CLUSTER_PARTIAL_READ (5921L)
value ERROR_CLUSTER_PARTIAL_SEND (5914L)
value ERROR_CLUSTER_PARTIAL_WRITE (5922L)
value ERROR_CLUSTER_POISONED (5907L)
value ERROR_CLUSTER_PROPERTY_DATA_TYPE_MISMATCH (5895L)
value ERROR_CLUSTER_QUORUMLOG_NOT_FOUND (5891L)
value ERROR_CLUSTER_REGISTRY_INVALID_FUNCTION (5915L)
value ERROR_CLUSTER_RESNAME_NOT_FOUND (5080L)
value ERROR_CLUSTER_RESOURCES_MUST_BE_ONLINE_ON_THE_SAME_NODE (5933L)
value ERROR_CLUSTER_RESOURCE_CONFIGURATION_ERROR (5943L)
value ERROR_CLUSTER_RESOURCE_CONTAINS_UNSUPPORTED_DIFF_AREA_FOR_SHARED_VOLUMES (5969L)
value ERROR_CLUSTER_RESOURCE_DOES_NOT_SUPPORT_UNMONITORED (5982L)
value ERROR_CLUSTER_RESOURCE_IS_IN_MAINTENANCE_MODE (5970L)
value ERROR_CLUSTER_RESOURCE_IS_REPLICATED (5983L)
value ERROR_CLUSTER_RESOURCE_IS_REPLICA_VIRTUAL_MACHINE (5972L)
value ERROR_CLUSTER_RESOURCE_LOCKED_STATUS (5960L)
value ERROR_CLUSTER_RESOURCE_NOT_MONITORED (5981L)
value ERROR_CLUSTER_RESOURCE_PROVIDER_FAILED (5942L)
value ERROR_CLUSTER_RESOURCE_TYPE_BUSY (5909L)
value ERROR_CLUSTER_RESOURCE_TYPE_NOT_FOUND (5078L)
value ERROR_CLUSTER_RESOURCE_VETOED_CALL (5955L)
value ERROR_CLUSTER_RESOURCE_VETOED_MOVE_INCOMPATIBLE_NODES (5953L)
value ERROR_CLUSTER_RESOURCE_VETOED_MOVE_NOT_ENOUGH_RESOURCES_ON_DESTINATION (5957L)
value ERROR_CLUSTER_RESOURCE_VETOED_MOVE_NOT_ENOUGH_RESOURCES_ON_SOURCE (5958L)
value ERROR_CLUSTER_RESTYPE_NOT_SUPPORTED (5079L)
value ERROR_CLUSTER_RHS_FAILED_INITIALIZATION (5931L)
value ERROR_CLUSTER_SHARED_VOLUMES_IN_USE (5947L)
value ERROR_CLUSTER_SHARED_VOLUME_FAILOVER_NOT_ALLOWED (5961L)
value ERROR_CLUSTER_SHARED_VOLUME_NOT_REDIRECTED (5967L)
value ERROR_CLUSTER_SHARED_VOLUME_REDIRECTED (5966L)
value ERROR_CLUSTER_SHUTTING_DOWN (5022L)
value ERROR_CLUSTER_SINGLETON_RESOURCE (5940L)
value ERROR_CLUSTER_SPACE_DEGRADED (5987L)
value ERROR_CLUSTER_SYSTEM_CONFIG_CHANGED (5077L)
value ERROR_CLUSTER_TOKEN_DELEGATION_NOT_SUPPORTED (5988L)
value ERROR_CLUSTER_TOO_MANY_NODES (5935L)
value ERROR_CLUSTER_UPGRADE_FIX_QUORUM_NOT_SUPPORTED (5974L)
value ERROR_CLUSTER_UPGRADE_INCOMPATIBLE_VERSIONS (5973L)
value ERROR_CLUSTER_UPGRADE_INCOMPLETE (5977L)
value ERROR_CLUSTER_UPGRADE_IN_PROGRESS (5976L)
value ERROR_CLUSTER_UPGRADE_RESTART_REQUIRED (5975L)
value ERROR_CLUSTER_USE_SHARED_VOLUMES_API (5948L)
value ERROR_CLUSTER_WATCHDOG_TERMINATING (5952L)
value ERROR_CLUSTER_WRONG_OS_VERSION (5899L)
value ERROR_COLORSPACE_MISMATCH (2021L)
value ERROR_COMMITMENT_LIMIT (1455L)
value ERROR_COMMITMENT_MINIMUM (635L)
value ERROR_COMPRESSED_FILE_NOT_SUPPORTED (335L)
value ERROR_COMPRESSION_DISABLED (769L)
value ERROR_COMPRESSION_NOT_ALLOWED_IN_TRANSACTION (6850L)
value ERROR_COMPRESSION_NOT_BENEFICIAL (344L)
value ERROR_COM_TASK_STOP_PENDING (15501L)
value ERROR_CONNECTED_OTHER_PASSWORD (2108L)
value ERROR_CONNECTED_OTHER_PASSWORD_DEFAULT (2109L)
value ERROR_CONNECTION_ABORTED (1236L)
value ERROR_CONNECTION_ACTIVE (1230L)
value ERROR_CONNECTION_COUNT_LIMIT (1238L)
value ERROR_CONNECTION_INVALID (1229L)
value ERROR_CONNECTION_REFUSED (1225L)
value ERROR_CONNECTION_UNAVAIL (1201L)
value ERROR_CONTAINER_ASSIGNED (1504L)
value ERROR_CONTENT_BLOCKED (1296L)
value ERROR_CONTEXT_EXPIRED (1931L)
value ERROR_CONTINUE (1246L)
value ERROR_CONTROLLING_IEPORT (4329L)
value ERROR_CONTROL_C_EXIT (572L)
value ERROR_CONTROL_ID_NOT_FOUND (1421L)
value ERROR_CONVERT_TO_LARGE (600L)
value ERROR_CORE_DRIVER_PACKAGE_NOT_FOUND (3016L)
value ERROR_CORE_RESOURCE (5026L)
value ERROR_CORRUPT_LOG_CLEARED (798L)
value ERROR_CORRUPT_LOG_CORRUPTED (795L)
value ERROR_CORRUPT_LOG_DELETED_FULL (797L)
value ERROR_CORRUPT_LOG_OVERFULL (794L)
value ERROR_CORRUPT_LOG_UNAVAILABLE (796L)
value ERROR_CORRUPT_SYSTEM_FILE (634L)
value ERROR_COULD_NOT_INTERPRET (552L)
value ERROR_COULD_NOT_RESIZE_LOG (6629L)
value ERROR_COUNTER_TIMEOUT (1121L)
value ERROR_CPU_SET_INVALID (813L)
value ERROR_CRASH_DUMP (753L)
value ERROR_CRC (23L)
value ERROR_CREATE_FAILED (1631L)
value ERROR_CRM_PROTOCOL_ALREADY_EXISTS (6710L)
value ERROR_CRM_PROTOCOL_NOT_FOUND (6712L)
value ERROR_CROSS_PARTITION_VIOLATION (1661L)
value ERROR_CSCSHARE_OFFLINE (1262L)
value ERROR_CSV_VOLUME_NOT_LOCAL (5951L)
value ERROR_CS_ENCRYPTION_EXISTING_ENCRYPTED_FILE (6019L)
value ERROR_CS_ENCRYPTION_FILE_NOT_CSE (6021L)
value ERROR_CS_ENCRYPTION_INVALID_SERVER_RESPONSE (6017L)
value ERROR_CS_ENCRYPTION_NEW_ENCRYPTED_FILE (6020L)
value ERROR_CS_ENCRYPTION_UNSUPPORTED_SERVER (6018L)
value ERROR_CTX_ACCOUNT_RESTRICTION (7064L)
value ERROR_CTX_BAD_VIDEO_MODE (7025L)
value ERROR_CTX_CANNOT_MAKE_EVENTLOG_ENTRY (7005L)
value ERROR_CTX_CDM_CONNECT (7066L)
value ERROR_CTX_CDM_DISCONNECT (7067L)
value ERROR_CTX_CLIENT_LICENSE_IN_USE (7052L)
value ERROR_CTX_CLIENT_LICENSE_NOT_SET (7053L)
value ERROR_CTX_CLIENT_QUERY_TIMEOUT (7040L)
value ERROR_CTX_CLOSE_PENDING (7007L)
value ERROR_CTX_CONSOLE_CONNECT (7042L)
value ERROR_CTX_CONSOLE_DISCONNECT (7041L)
value ERROR_CTX_ENCRYPTION_LEVEL_REQUIRED (7061L)
value ERROR_CTX_GRAPHICS_INVALID (7035L)
value ERROR_CTX_INVALID_MODEMNAME (7010L)
value ERROR_CTX_INVALID_PD (7002L)
value ERROR_CTX_INVALID_WD (7049L)
value ERROR_CTX_LICENSE_CLIENT_INVALID (7055L)
value ERROR_CTX_LICENSE_EXPIRED (7056L)
value ERROR_CTX_LICENSE_NOT_AVAILABLE (7054L)
value ERROR_CTX_LOGON_DISABLED (7037L)
value ERROR_CTX_MODEM_INF_NOT_FOUND (7009L)
value ERROR_CTX_MODEM_RESPONSE_BUSY (7015L)
value ERROR_CTX_MODEM_RESPONSE_ERROR (7011L)
value ERROR_CTX_MODEM_RESPONSE_NO_CARRIER (7013L)
value ERROR_CTX_MODEM_RESPONSE_NO_DIALTONE (7014L)
value ERROR_CTX_MODEM_RESPONSE_TIMEOUT (7012L)
value ERROR_CTX_MODEM_RESPONSE_VOICE (7016L)
value ERROR_CTX_NOT_CONSOLE (7038L)
value ERROR_CTX_NO_FORCE_LOGOFF (7063L)
value ERROR_CTX_NO_OUTBUF (7008L)
value ERROR_CTX_PD_NOT_FOUND (7003L)
value ERROR_CTX_SECURITY_LAYER_ERROR (7068L)
value ERROR_CTX_SERVICE_NAME_COLLISION (7006L)
value ERROR_CTX_SESSION_IN_USE (7062L)
value ERROR_CTX_SHADOW_DENIED (7044L)
value ERROR_CTX_SHADOW_DISABLED (7051L)
value ERROR_CTX_SHADOW_ENDED_BY_MODE_CHANGE (7058L)
value ERROR_CTX_SHADOW_INVALID (7050L)
value ERROR_CTX_SHADOW_NOT_RUNNING (7057L)
value ERROR_CTX_TD_ERROR (7017L)
value ERROR_CTX_WD_NOT_FOUND (7004L)
value ERROR_CTX_WINSTATIONS_DISABLED (7060L)
value ERROR_CTX_WINSTATION_ACCESS_DENIED (7045L)
value ERROR_CTX_WINSTATION_ALREADY_EXISTS (7023L)
value ERROR_CTX_WINSTATION_BUSY (7024L)
value ERROR_CTX_WINSTATION_NAME_INVALID (7001L)
value ERROR_CTX_WINSTATION_NOT_FOUND (7022L)
value ERROR_CURRENT_DIRECTORY (16L)
value ERROR_CURRENT_DOMAIN_NOT_ALLOWED (1399L)
value ERROR_CURRENT_TRANSACTION_NOT_VALID (6714L)
value ERROR_DATABASE_BACKUP_CORRUPT (5087L)
value ERROR_DATABASE_DOES_NOT_EXIST (1065L)
value ERROR_DATABASE_FAILURE (4313L)
value ERROR_DATABASE_FULL (4314L)
value ERROR_DATATYPE_MISMATCH (1629L)
value ERROR_DATA_CHECKSUM_ERROR (323L)
value ERROR_DATA_LOST_REPAIR (6843L)
value ERROR_DATA_NOT_ACCEPTED (592L)
value ERROR_DAX_MAPPING_EXISTS (361L)
value ERROR_DBG_COMMAND_EXCEPTION (697L)
value ERROR_DBG_CONTINUE (767L)
value ERROR_DBG_CONTROL_BREAK (696L)
value ERROR_DBG_CONTROL_C (693L)
value ERROR_DBG_EXCEPTION_HANDLED (766L)
value ERROR_DBG_EXCEPTION_NOT_HANDLED (688L)
value ERROR_DBG_PRINTEXCEPTION_C (694L)
value ERROR_DBG_REPLY_LATER (689L)
value ERROR_DBG_RIPEXCEPTION (695L)
value ERROR_DBG_TERMINATE_PROCESS (692L)
value ERROR_DBG_TERMINATE_THREAD (691L)
value ERROR_DBG_UNABLE_TO_PROVIDE_HANDLE (690L)
value ERROR_DC_NOT_FOUND (1425L)
value ERROR_DDE_FAIL (1156L)
value ERROR_DEBUGGER_INACTIVE (1284L)
value ERROR_DEBUG_ATTACH_FAILED (590L)
value ERROR_DECRYPTION_FAILED (6001L)
value ERROR_DELAY_LOAD_FAILED (1285L)
value ERROR_DELETE_PENDING (303L)
value ERROR_DELETING_EXISTING_APPLICATIONDATA_STORE_FAILED (15621L)
value ERROR_DELETING_ICM_XFORM (2019L)
value ERROR_DEPENDENCY_ALREADY_EXISTS (5003L)
value ERROR_DEPENDENCY_NOT_ALLOWED (5069L)
value ERROR_DEPENDENCY_NOT_FOUND (5002L)
value ERROR_DEPENDENCY_TREE_TOO_COMPLEX (5929L)
value ERROR_DEPENDENT_RESOURCE_EXISTS (5001L)
value ERROR_DEPENDENT_RESOURCE_PROPERTY_CONFLICT (5924L)
value ERROR_DEPENDENT_SERVICES_RUNNING (1051L)
value ERROR_DEPLOYMENT_BLOCKED_BY_POLICY (15617L)
value ERROR_DEPLOYMENT_BLOCKED_BY_PROFILE_POLICY (15651L)
value ERROR_DEPLOYMENT_BLOCKED_BY_USER_LOG_OFF (15641L)
value ERROR_DEPLOYMENT_BLOCKED_BY_VOLUME_POLICY_MACHINE (15650L)
value ERROR_DEPLOYMENT_BLOCKED_BY_VOLUME_POLICY_PACKAGE (15649L)
value ERROR_DEPLOYMENT_FAILED_CONFLICTING_MUTABLE_PACKAGE_DIRECTORY (15652L)
value ERROR_DEPLOYMENT_OPTION_NOT_SUPPORTED (15645L)
value ERROR_DESTINATION_ELEMENT_FULL (1161L)
value ERROR_DESTROY_OBJECT_OF_OTHER_THREAD (1435L)
value ERROR_DEVICE_ALREADY_ATTACHED (548L)
value ERROR_DEVICE_ALREADY_REMEMBERED (1202L)
value ERROR_DEVICE_DOOR_OPEN (1166L)
value ERROR_DEVICE_ENUMERATION_ERROR (648L)
value ERROR_DEVICE_FEATURE_NOT_SUPPORTED (316L)
value ERROR_DEVICE_HARDWARE_ERROR (483L)
value ERROR_DEVICE_HINT_NAME_BUFFER_TOO_SMALL (355L)
value ERROR_DEVICE_IN_MAINTENANCE (359L)
value ERROR_DEVICE_IN_USE (2404L)
value ERROR_DEVICE_NOT_AVAILABLE (4319L)
value ERROR_DEVICE_NOT_CONNECTED (1167L)
value ERROR_DEVICE_NOT_PARTITIONED (1107L)
value ERROR_DEVICE_NO_RESOURCES (322L)
value ERROR_DEVICE_REINITIALIZATION_NEEDED (1164L)
value ERROR_DEVICE_REMOVED (1617L)
value ERROR_DEVICE_REQUIRES_CLEANING (1165L)
value ERROR_DEVICE_RESET_REQUIRED (507L)
value ERROR_DEVICE_SUPPORT_IN_PROGRESS (171L)
value ERROR_DEVICE_UNREACHABLE (321L)
value ERROR_DEV_NOT_EXIST (55L)
value ERROR_DEV_SIDELOAD_LIMIT_EXCEEDED (15633L)
value ERROR_DHCP_ADDRESS_CONFLICT (4100L)
value ERROR_DIFFERENT_PROFILE_RESOURCE_MANAGER_EXIST (15144L)
value ERROR_DIFFERENT_SERVICE_ACCOUNT (1079L)
value ERROR_DIFFERENT_VERSION_OF_PACKAGED_SERVICE_INSTALLED (15654L)
value ERROR_DIF_BINDING_API_NOT_FOUND (3199L)
value ERROR_DIF_IOCALLBACK_NOT_REPLACED (3190L)
value ERROR_DIF_LIVEDUMP_LIMIT_EXCEEDED (3191L)
value ERROR_DIF_VOLATILE_DRIVER_HOTPATCHED (3193L)
value ERROR_DIF_VOLATILE_DRIVER_IS_NOT_RUNNING (3195L)
value ERROR_DIF_VOLATILE_INVALID_INFO (3194L)
value ERROR_DIF_VOLATILE_NOT_ALLOWED (3198L)
value ERROR_DIF_VOLATILE_PLUGIN_CHANGE_NOT_ALLOWED (3197L)
value ERROR_DIF_VOLATILE_PLUGIN_IS_NOT_RUNNING (3196L)
value ERROR_DIF_VOLATILE_SECTION_NOT_LOCKED (3192L)
value ERROR_DIRECTORY (267L)
value ERROR_DIRECTORY_NOT_RM (6803L)
value ERROR_DIRECTORY_NOT_SUPPORTED (336L)
value ERROR_DIRECT_ACCESS_HANDLE (130L)
value ERROR_DIR_EFS_DISALLOWED (6010L)
value ERROR_DIR_NOT_EMPTY (145L)
value ERROR_DIR_NOT_ROOT (144L)
value ERROR_DISCARDED (157L)
value ERROR_DISK_CHANGE (107L)
value ERROR_DISK_CORRUPT (1393L)
value ERROR_DISK_FULL (112L)
value ERROR_DISK_NOT_CSV_CAPABLE (5964L)
value ERROR_DISK_OPERATION_FAILED (1127L)
value ERROR_DISK_QUOTA_EXCEEDED (1295L)
value ERROR_DISK_RECALIBRATE_FAILED (1126L)
value ERROR_DISK_REPAIR_DISABLED (780L)
value ERROR_DISK_REPAIR_REDIRECTED (792L)
value ERROR_DISK_REPAIR_UNSUCCESSFUL (793L)
value ERROR_DISK_RESET_FAILED (1128L)
value ERROR_DISK_RESOURCES_EXHAUSTED (314L)
value ERROR_DISK_TOO_FRAGMENTED (302L)
value ERROR_DLL_INIT_FAILED (1114L)
value ERROR_DLL_INIT_FAILED_LOGOFF (624L)
value ERROR_DLL_MIGHT_BE_INCOMPATIBLE (687L)
value ERROR_DLL_MIGHT_BE_INSECURE (686L)
value ERROR_DLL_NOT_FOUND (1157L)
value ERROR_DLP_POLICY_DENIES_OPERATION (446L)
value ERROR_DLP_POLICY_SILENTLY_FAIL (449L)
value ERROR_DLP_POLICY_WARNS_AGAINST_OPERATION (445L)
value ERROR_DOMAIN_CONTROLLER_EXISTS (1250L)
value ERROR_DOMAIN_CONTROLLER_NOT_FOUND (1908L)
value ERROR_DOMAIN_CTRLR_CONFIG_ERROR (581L)
value ERROR_DOMAIN_EXISTS (1356L)
value ERROR_DOMAIN_LIMIT_EXCEEDED (1357L)
value ERROR_DOMAIN_SID_SAME_AS_LOCAL_WORKSTATION (8644L)
value ERROR_DOMAIN_TRUST_INCONSISTENT (1810L)
value ERROR_DOWNGRADE_DETECTED (1265L)
value ERROR_DPL_NOT_SUPPORTED_FOR_USER (423L)
value ERROR_DRIVERS_LEAKING_LOCKED_PAGES (729L)
value ERROR_DRIVER_BLOCKED (1275L)
value ERROR_DRIVER_CANCEL_TIMEOUT (594L)
value ERROR_DRIVER_DATABASE_ERROR (652L)
value ERROR_DRIVER_FAILED_PRIOR_UNLOAD (654L)
value ERROR_DRIVER_FAILED_SLEEP (633L)
value ERROR_DRIVER_PROCESS_TERMINATED (1291L)
value ERROR_DRIVE_LOCKED (108L)
value ERROR_DRIVE_MEDIA_MISMATCH (4303L)
value ERROR_DS_ADD_REPLICA_INHIBITED (8302L)
value ERROR_DS_ADMIN_LIMIT_EXCEEDED (8228L)
value ERROR_DS_AFFECTS_MULTIPLE_DSAS (8249L)
value ERROR_DS_AG_CANT_HAVE_UNIVERSAL_MEMBER (8578L)
value ERROR_DS_ALIASED_OBJ_MISSING (8334L)
value ERROR_DS_ALIAS_DEREF_PROBLEM (8244L)
value ERROR_DS_ALIAS_POINTS_TO_ALIAS (8336L)
value ERROR_DS_ALIAS_PROBLEM (8241L)
value ERROR_DS_ATTRIBUTE_OR_VALUE_EXISTS (8205L)
value ERROR_DS_ATTRIBUTE_OWNED_BY_SAM (8346L)
value ERROR_DS_ATTRIBUTE_TYPE_UNDEFINED (8204L)
value ERROR_DS_ATT_ALREADY_EXISTS (8318L)
value ERROR_DS_ATT_IS_NOT_ON_OBJ (8310L)
value ERROR_DS_ATT_NOT_DEF_FOR_CLASS (8317L)
value ERROR_DS_ATT_NOT_DEF_IN_SCHEMA (8303L)
value ERROR_DS_ATT_SCHEMA_REQ_ID (8399L)
value ERROR_DS_ATT_SCHEMA_REQ_SYNTAX (8416L)
value ERROR_DS_ATT_VAL_ALREADY_EXISTS (8323L)
value ERROR_DS_AUDIT_FAILURE (8625L)
value ERROR_DS_AUTHORIZATION_FAILED (8599L)
value ERROR_DS_AUTH_METHOD_NOT_SUPPORTED (8231L)
value ERROR_DS_AUTH_UNKNOWN (8234L)
value ERROR_DS_AUX_CLS_TEST_FAIL (8389L)
value ERROR_DS_BACKLINK_WITHOUT_LINK (8482L)
value ERROR_DS_BAD_ATT_SCHEMA_SYNTAX (8400L)
value ERROR_DS_BAD_HIERARCHY_FILE (8425L)
value ERROR_DS_BAD_INSTANCE_TYPE (8313L)
value ERROR_DS_BAD_NAME_SYNTAX (8335L)
value ERROR_DS_BAD_RDN_ATT_ID_SYNTAX (8392L)
value ERROR_DS_BUILD_HIERARCHY_TABLE_FAILED (8426L)
value ERROR_DS_BUSY (8206L)
value ERROR_DS_CANT_ACCESS_REMOTE_PART_OF_AD (8585L)
value ERROR_DS_CANT_ADD_ATT_VALUES (8320L)
value ERROR_DS_CANT_ADD_SYSTEM_ONLY (8358L)
value ERROR_DS_CANT_ADD_TO_GC (8550L)
value ERROR_DS_CANT_CACHE_ATT (8401L)
value ERROR_DS_CANT_CACHE_CLASS (8402L)
value ERROR_DS_CANT_CREATE_IN_NONDOMAIN_NC (8553L)
value ERROR_DS_CANT_CREATE_UNDER_SCHEMA (8510L)
value ERROR_DS_CANT_DELETE (8398L)
value ERROR_DS_CANT_DELETE_DSA_OBJ (8340L)
value ERROR_DS_CANT_DEL_MASTER_CROSSREF (8375L)
value ERROR_DS_CANT_DEMOTE_WITH_WRITEABLE_NC (8604L)
value ERROR_DS_CANT_DEREF_ALIAS (8337L)
value ERROR_DS_CANT_DERIVE_SPN_FOR_DELETED_DOMAIN (8603L)
value ERROR_DS_CANT_DERIVE_SPN_WITHOUT_SERVER_REF (8589L)
value ERROR_DS_CANT_FIND_DC_FOR_SRC_DOMAIN (8537L)
value ERROR_DS_CANT_FIND_DSA_OBJ (8419L)
value ERROR_DS_CANT_FIND_EXPECTED_NC (8420L)
value ERROR_DS_CANT_FIND_NC_IN_CACHE (8421L)
value ERROR_DS_CANT_MIX_MASTER_AND_REPS (8331L)
value ERROR_DS_CANT_MOD_OBJ_CLASS (8215L)
value ERROR_DS_CANT_MOD_PRIMARYGROUPID (8506L)
value ERROR_DS_CANT_MOD_SYSTEM_ONLY (8369L)
value ERROR_DS_CANT_MOVE_ACCOUNT_GROUP (8498L)
value ERROR_DS_CANT_MOVE_APP_BASIC_GROUP (8608L)
value ERROR_DS_CANT_MOVE_APP_QUERY_GROUP (8609L)
value ERROR_DS_CANT_MOVE_DELETED_OBJECT (8489L)
value ERROR_DS_CANT_MOVE_RESOURCE_GROUP (8499L)
value ERROR_DS_CANT_ON_NON_LEAF (8213L)
value ERROR_DS_CANT_ON_RDN (8214L)
value ERROR_DS_CANT_REMOVE_ATT_CACHE (8403L)
value ERROR_DS_CANT_REMOVE_CLASS_CACHE (8404L)
value ERROR_DS_CANT_REM_MISSING_ATT (8324L)
value ERROR_DS_CANT_REM_MISSING_ATT_VAL (8325L)
value ERROR_DS_CANT_REPLACE_HIDDEN_REC (8424L)
value ERROR_DS_CANT_RETRIEVE_ATTS (8481L)
value ERROR_DS_CANT_RETRIEVE_CHILD (8422L)
value ERROR_DS_CANT_RETRIEVE_DN (8405L)
value ERROR_DS_CANT_RETRIEVE_INSTANCE (8407L)
value ERROR_DS_CANT_RETRIEVE_SD (8526L)
value ERROR_DS_CANT_START (8531L)
value ERROR_DS_CANT_TREE_DELETE_CRITICAL_OBJ (8560L)
value ERROR_DS_CANT_WITH_ACCT_GROUP_MEMBERSHPS (8493L)
value ERROR_DS_CHILDREN_EXIST (8332L)
value ERROR_DS_CLASS_MUST_BE_CONCRETE (8359L)
value ERROR_DS_CLASS_NOT_DSA (8343L)
value ERROR_DS_CLIENT_LOOP (8259L)
value ERROR_DS_CODE_INCONSISTENCY (8408L)
value ERROR_DS_COMPARE_FALSE (8229L)
value ERROR_DS_COMPARE_TRUE (8230L)
value ERROR_DS_CONFIDENTIALITY_REQUIRED (8237L)
value ERROR_DS_CONFIG_PARAM_MISSING (8427L)
value ERROR_DS_CONSTRAINT_VIOLATION (8239L)
value ERROR_DS_CONSTRUCTED_ATT_MOD (8475L)
value ERROR_DS_CONTROL_NOT_FOUND (8258L)
value ERROR_DS_COULDNT_CONTACT_FSMO (8367L)
value ERROR_DS_COULDNT_IDENTIFY_OBJECTS_FOR_TREE_DELETE (8503L)
value ERROR_DS_COULDNT_LOCK_TREE_FOR_DELETE (8502L)
value ERROR_DS_COULDNT_UPDATE_SPNS (8525L)
value ERROR_DS_COUNTING_AB_INDICES_FAILED (8428L)
value ERROR_DS_CROSS_DOMAIN_CLEANUP_REQD (8491L)
value ERROR_DS_CROSS_DOM_MOVE_ERROR (8216L)
value ERROR_DS_CROSS_NC_DN_RENAME (8368L)
value ERROR_DS_CROSS_REF_BUSY (8602L)
value ERROR_DS_CROSS_REF_EXISTS (8374L)
value ERROR_DS_CR_IMPOSSIBLE_TO_VALIDATE (8495L)
value ERROR_DS_DATABASE_ERROR (8409L)
value ERROR_DS_DECODING_ERROR (8253L)
value ERROR_DS_DESTINATION_AUDITING_NOT_ENABLED (8536L)
value ERROR_DS_DESTINATION_DOMAIN_NOT_IN_FOREST (8535L)
value ERROR_DS_DIFFERENT_REPL_EPOCHS (8593L)
value ERROR_DS_DISALLOWED_IN_SYSTEM_CONTAINER (8615L)
value ERROR_DS_DISALLOWED_NC_REDIRECT (8640L)
value ERROR_DS_DNS_LOOKUP_FAILURE (8524L)
value ERROR_DS_DOMAIN_NAME_EXISTS_IN_FOREST (8634L)
value ERROR_DS_DOMAIN_RENAME_IN_PROGRESS (8612L)
value ERROR_DS_DOMAIN_VERSION_TOO_HIGH (8564L)
value ERROR_DS_DOMAIN_VERSION_TOO_LOW (8566L)
value ERROR_DS_DRA_ABANDON_SYNC (8462L)
value ERROR_DS_DRA_ACCESS_DENIED (8453L)
value ERROR_DS_DRA_BAD_DN (8439L)
value ERROR_DS_DRA_BAD_INSTANCE_TYPE (8445L)
value ERROR_DS_DRA_BAD_NC (8440L)
value ERROR_DS_DRA_BUSY (8438L)
value ERROR_DS_DRA_CONNECTION_FAILED (8444L)
value ERROR_DS_DRA_CORRUPT_UTD_VECTOR (8629L)
value ERROR_DS_DRA_DB_ERROR (8451L)
value ERROR_DS_DRA_DN_EXISTS (8441L)
value ERROR_DS_DRA_EARLIER_SCHEMA_CONFLICT (8544L)
value ERROR_DS_DRA_EXTN_CONNECTION_FAILED (8466L)
value ERROR_DS_DRA_GENERIC (8436L)
value ERROR_DS_DRA_INCOMPATIBLE_PARTIAL_SET (8464L)
value ERROR_DS_DRA_INCONSISTENT_DIT (8443L)
value ERROR_DS_DRA_INTERNAL_ERROR (8442L)
value ERROR_DS_DRA_INVALID_PARAMETER (8437L)
value ERROR_DS_DRA_MAIL_PROBLEM (8447L)
value ERROR_DS_DRA_MISSING_KRBTGT_SECRET (8633L)
value ERROR_DS_DRA_MISSING_PARENT (8460L)
value ERROR_DS_DRA_NAME_COLLISION (8458L)
value ERROR_DS_DRA_NOT_SUPPORTED (8454L)
value ERROR_DS_DRA_NO_REPLICA (8452L)
value ERROR_DS_DRA_OBJ_IS_REP_SOURCE (8450L)
value ERROR_DS_DRA_OBJ_NC_MISMATCH (8545L)
value ERROR_DS_DRA_OUT_OF_MEM (8446L)
value ERROR_DS_DRA_OUT_SCHEDULE_WINDOW (8617L)
value ERROR_DS_DRA_PREEMPTED (8461L)
value ERROR_DS_DRA_RECYCLED_TARGET (8639L)
value ERROR_DS_DRA_REF_ALREADY_EXISTS (8448L)
value ERROR_DS_DRA_REF_NOT_FOUND (8449L)
value ERROR_DS_DRA_REPL_PENDING (8477L)
value ERROR_DS_DRA_RPC_CANCELLED (8455L)
value ERROR_DS_DRA_SCHEMA_CONFLICT (8543L)
value ERROR_DS_DRA_SCHEMA_INFO_SHIP (8542L)
value ERROR_DS_DRA_SCHEMA_MISMATCH (8418L)
value ERROR_DS_DRA_SECRETS_DENIED (8630L)
value ERROR_DS_DRA_SHUTDOWN (8463L)
value ERROR_DS_DRA_SINK_DISABLED (8457L)
value ERROR_DS_DRA_SOURCE_DISABLED (8456L)
value ERROR_DS_DRA_SOURCE_IS_PARTIAL_REPLICA (8465L)
value ERROR_DS_DRA_SOURCE_REINSTALLED (8459L)
value ERROR_DS_DRS_EXTENSIONS_CHANGED (8594L)
value ERROR_DS_DSA_MUST_BE_INT_MASTER (8342L)
value ERROR_DS_DST_DOMAIN_NOT_NATIVE (8496L)
value ERROR_DS_DST_NC_MISMATCH (8486L)
value ERROR_DS_DS_REQUIRED (8478L)
value ERROR_DS_DUPLICATE_ID_FOUND (8605L)
value ERROR_DS_DUP_LDAP_DISPLAY_NAME (8382L)
value ERROR_DS_DUP_LINK_ID (8468L)
value ERROR_DS_DUP_MAPI_ID (8380L)
value ERROR_DS_DUP_MSDS_INTID (8597L)
value ERROR_DS_DUP_OID (8379L)
value ERROR_DS_DUP_RDN (8378L)
value ERROR_DS_DUP_SCHEMA_ID_GUID (8381L)
value ERROR_DS_ENCODING_ERROR (8252L)
value ERROR_DS_EPOCH_MISMATCH (8483L)
value ERROR_DS_EXISTING_AD_CHILD_NC (8613L)
value ERROR_DS_EXISTS_IN_AUX_CLS (8393L)
value ERROR_DS_EXISTS_IN_MAY_HAVE (8386L)
value ERROR_DS_EXISTS_IN_MUST_HAVE (8385L)
value ERROR_DS_EXISTS_IN_POSS_SUP (8395L)
value ERROR_DS_EXISTS_IN_RDNATTID (8598L)
value ERROR_DS_EXISTS_IN_SUB_CLS (8394L)
value ERROR_DS_FILTER_UNKNOWN (8254L)
value ERROR_DS_FILTER_USES_CONTRUCTED_ATTRS (8555L)
value ERROR_DS_FLAT_NAME_EXISTS_IN_FOREST (8635L)
value ERROR_DS_FOREST_VERSION_TOO_HIGH (8563L)
value ERROR_DS_FOREST_VERSION_TOO_LOW (8565L)
value ERROR_DS_GCVERIFY_ERROR (8417L)
value ERROR_DS_GC_NOT_AVAILABLE (8217L)
value ERROR_DS_GC_REQUIRED (8547L)
value ERROR_DS_GENERIC_ERROR (8341L)
value ERROR_DS_GLOBAL_CANT_HAVE_CROSSDOMAIN_MEMBER (8519L)
value ERROR_DS_GLOBAL_CANT_HAVE_LOCAL_MEMBER (8516L)
value ERROR_DS_GLOBAL_CANT_HAVE_UNIVERSAL_MEMBER (8517L)
value ERROR_DS_GOVERNSID_MISSING (8410L)
value ERROR_DS_GROUP_CONVERSION_ERROR (8607L)
value ERROR_DS_HAVE_PRIMARY_MEMBERS (8521L)
value ERROR_DS_HIERARCHY_TABLE_MALLOC_FAILED (8429L)
value ERROR_DS_HIERARCHY_TABLE_TOO_DEEP (8628L)
value ERROR_DS_HIGH_ADLDS_FFL (8641L)
value ERROR_DS_HIGH_DSA_VERSION (8642L)
value ERROR_DS_ILLEGAL_BASE_SCHEMA_MOD (8507L)
value ERROR_DS_ILLEGAL_MOD_OPERATION (8311L)
value ERROR_DS_ILLEGAL_SUPERIOR (8345L)
value ERROR_DS_ILLEGAL_XDOM_MOVE_OPERATION (8492L)
value ERROR_DS_INAPPROPRIATE_AUTH (8233L)
value ERROR_DS_INAPPROPRIATE_MATCHING (8238L)
value ERROR_DS_INCOMPATIBLE_CONTROLS_USED (8574L)
value ERROR_DS_INCOMPATIBLE_VERSION (8567L)
value ERROR_DS_INCORRECT_ROLE_OWNER (8210L)
value ERROR_DS_INIT_FAILURE (8532L)
value ERROR_DS_INIT_FAILURE_CONSOLE (8561L)
value ERROR_DS_INSTALL_NO_SCH_VERSION_IN_INIFILE (8512L)
value ERROR_DS_INSTALL_NO_SRC_SCH_VERSION (8511L)
value ERROR_DS_INSTALL_SCHEMA_MISMATCH (8467L)
value ERROR_DS_INSUFFICIENT_ATTR_TO_CREATE_OBJECT (8606L)
value ERROR_DS_INSUFF_ACCESS_RIGHTS (8344L)
value ERROR_DS_INTERNAL_FAILURE (8430L)
value ERROR_DS_INVALID_ATTRIBUTE_SYNTAX (8203L)
value ERROR_DS_INVALID_DMD (8360L)
value ERROR_DS_INVALID_DN_SYNTAX (8242L)
value ERROR_DS_INVALID_GROUP_TYPE (8513L)
value ERROR_DS_INVALID_LDAP_DISPLAY_NAME (8479L)
value ERROR_DS_INVALID_NAME_FOR_SPN (8554L)
value ERROR_DS_INVALID_ROLE_OWNER (8366L)
value ERROR_DS_INVALID_SCRIPT (8600L)
value ERROR_DS_INVALID_SEARCH_FLAG (8500L)
value ERROR_DS_INVALID_SEARCH_FLAG_SUBTREE (8626L)
value ERROR_DS_INVALID_SEARCH_FLAG_TUPLE (8627L)
value ERROR_DS_IS_LEAF (8243L)
value ERROR_DS_KEY_NOT_UNIQUE (8527L)
value ERROR_DS_LDAP_SEND_QUEUE_FULL (8616L)
value ERROR_DS_LINK_ID_NOT_AVAILABLE (8577L)
value ERROR_DS_LOCAL_CANT_HAVE_CROSSDOMAIN_LOCAL_MEMBER (8520L)
value ERROR_DS_LOCAL_ERROR (8251L)
value ERROR_DS_LOCAL_MEMBER_OF_LOCAL_ONLY (8548L)
value ERROR_DS_LOOP_DETECT (8246L)
value ERROR_DS_LOW_ADLDS_FFL (8643L)
value ERROR_DS_LOW_DSA_VERSION (8568L)
value ERROR_DS_MACHINE_ACCOUNT_QUOTA_EXCEEDED (8557L)
value ERROR_DS_MAPI_ID_NOT_AVAILABLE (8632L)
value ERROR_DS_MASTERDSA_REQUIRED (8314L)
value ERROR_DS_MAX_OBJ_SIZE_EXCEEDED (8304L)
value ERROR_DS_MEMBERSHIP_EVALUATED_LOCALLY (8201L)
value ERROR_DS_MISSING_EXPECTED_ATT (8411L)
value ERROR_DS_MISSING_FOREST_TRUST (8649L)
value ERROR_DS_MISSING_FSMO_SETTINGS (8434L)
value ERROR_DS_MISSING_INFRASTRUCTURE_CONTAINER (8497L)
value ERROR_DS_MISSING_REQUIRED_ATT (8316L)
value ERROR_DS_MISSING_SUPREF (8406L)
value ERROR_DS_MODIFYDN_DISALLOWED_BY_FLAG (8581L)
value ERROR_DS_MODIFYDN_DISALLOWED_BY_INSTANCE_TYPE (8579L)
value ERROR_DS_MODIFYDN_WRONG_GRANDPARENT (8582L)
value ERROR_DS_MUST_BE_RUN_ON_DST_DC (8558L)
value ERROR_DS_NAME_ERROR_DOMAIN_ONLY (8473L)
value ERROR_DS_NAME_ERROR_NOT_FOUND (8470L)
value ERROR_DS_NAME_ERROR_NOT_UNIQUE (8471L)
value ERROR_DS_NAME_ERROR_NO_MAPPING (8472L)
value ERROR_DS_NAME_ERROR_NO_SYNTACTICAL_MAPPING (8474L)
value ERROR_DS_NAME_ERROR_RESOLVING (8469L)
value ERROR_DS_NAME_ERROR_TRUST_REFERRAL (8583L)
value ERROR_DS_NAME_NOT_UNIQUE (8571L)
value ERROR_DS_NAME_REFERENCE_INVALID (8373L)
value ERROR_DS_NAME_TOO_LONG (8348L)
value ERROR_DS_NAME_TOO_MANY_PARTS (8347L)
value ERROR_DS_NAME_TYPE_UNKNOWN (8351L)
value ERROR_DS_NAME_UNPARSEABLE (8350L)
value ERROR_DS_NAME_VALUE_TOO_LONG (8349L)
value ERROR_DS_NAMING_MASTER_GC (8523L)
value ERROR_DS_NAMING_VIOLATION (8247L)
value ERROR_DS_NCNAME_MISSING_CR_REF (8412L)
value ERROR_DS_NCNAME_MUST_BE_NC (8357L)
value ERROR_DS_NC_MUST_HAVE_NC_PARENT (8494L)
value ERROR_DS_NC_STILL_HAS_DSAS (8546L)
value ERROR_DS_NONEXISTENT_MAY_HAVE (8387L)
value ERROR_DS_NONEXISTENT_MUST_HAVE (8388L)
value ERROR_DS_NONEXISTENT_POSS_SUP (8390L)
value ERROR_DS_NONSAFE_SCHEMA_CHANGE (8508L)
value ERROR_DS_NON_ASQ_SEARCH (8624L)
value ERROR_DS_NON_BASE_SEARCH (8480L)
value ERROR_DS_NOTIFY_FILTER_TOO_COMPLEX (8377L)
value ERROR_DS_NOT_AN_OBJECT (8352L)
value ERROR_DS_NOT_AUTHORITIVE_FOR_DST_NC (8487L)
value ERROR_DS_NOT_CLOSEST (8588L)
value ERROR_DS_NOT_INSTALLED (8200L)
value ERROR_DS_NOT_ON_BACKLINK (8362L)
value ERROR_DS_NOT_SUPPORTED (8256L)
value ERROR_DS_NOT_SUPPORTED_SORT_ORDER (8570L)
value ERROR_DS_NO_ATTRIBUTE_OR_VALUE (8202L)
value ERROR_DS_NO_BEHAVIOR_VERSION_IN_MIXEDDOMAIN (8569L)
value ERROR_DS_NO_CHAINED_EVAL (8328L)
value ERROR_DS_NO_CHAINING (8327L)
value ERROR_DS_NO_CHECKPOINT_WITH_PDC (8551L)
value ERROR_DS_NO_CROSSREF_FOR_NC (8363L)
value ERROR_DS_NO_DELETED_NAME (8355L)
value ERROR_DS_NO_FPO_IN_UNIVERSAL_GROUPS (8549L)
value ERROR_DS_NO_MORE_RIDS (8209L)
value ERROR_DS_NO_MSDS_INTID (8596L)
value ERROR_DS_NO_NEST_GLOBALGROUP_IN_MIXEDDOMAIN (8514L)
value ERROR_DS_NO_NEST_LOCALGROUP_IN_MIXEDDOMAIN (8515L)
value ERROR_DS_NO_NTDSA_OBJECT (8623L)
value ERROR_DS_NO_OBJECT_MOVE_IN_SCHEMA_NC (8580L)
value ERROR_DS_NO_PARENT_OBJECT (8329L)
value ERROR_DS_NO_PKT_PRIVACY_ON_CONNECTION (8533L)
value ERROR_DS_NO_RDN_DEFINED_IN_SCHEMA (8306L)
value ERROR_DS_NO_REF_DOMAIN (8575L)
value ERROR_DS_NO_REQUESTED_ATTS_FOUND (8308L)
value ERROR_DS_NO_RESULTS_RETURNED (8257L)
value ERROR_DS_NO_RIDS_ALLOCATED (8208L)
value ERROR_DS_NO_SERVER_OBJECT (8622L)
value ERROR_DS_NO_SUCH_OBJECT (8240L)
value ERROR_DS_NO_TREE_DELETE_ABOVE_NC (8501L)
value ERROR_DS_NTDSCRIPT_PROCESS_ERROR (8592L)
value ERROR_DS_NTDSCRIPT_SYNTAX_ERROR (8591L)
value ERROR_DS_OBJECT_BEING_REMOVED (8339L)
value ERROR_DS_OBJECT_CLASS_REQUIRED (8315L)
value ERROR_DS_OBJECT_RESULTS_TOO_LARGE (8248L)
value ERROR_DS_OBJ_CLASS_NOT_DEFINED (8371L)
value ERROR_DS_OBJ_CLASS_NOT_SUBCLASS (8372L)
value ERROR_DS_OBJ_CLASS_VIOLATION (8212L)
value ERROR_DS_OBJ_GUID_EXISTS (8361L)
value ERROR_DS_OBJ_NOT_FOUND (8333L)
value ERROR_DS_OBJ_STRING_NAME_EXISTS (8305L)
value ERROR_DS_OBJ_TOO_LARGE (8312L)
value ERROR_DS_OFFSET_RANGE_ERROR (8262L)
value ERROR_DS_OID_MAPPED_GROUP_CANT_HAVE_MEMBERS (8637L)
value ERROR_DS_OID_NOT_FOUND (8638L)
value ERROR_DS_OPERATIONS_ERROR (8224L)
value ERROR_DS_OUT_OF_SCOPE (8338L)
value ERROR_DS_OUT_OF_VERSION_STORE (8573L)
value ERROR_DS_PARAM_ERROR (8255L)
value ERROR_DS_PARENT_IS_AN_ALIAS (8330L)
value ERROR_DS_PDC_OPERATION_IN_PROGRESS (8490L)
value ERROR_DS_PER_ATTRIBUTE_AUTHZ_FAILED_DURING_ADD (8652L)
value ERROR_DS_POLICY_NOT_KNOWN (8618L)
value ERROR_DS_PROTOCOL_ERROR (8225L)
value ERROR_DS_RANGE_CONSTRAINT (8322L)
value ERROR_DS_RDN_DOESNT_MATCH_SCHEMA (8307L)
value ERROR_DS_RECALCSCHEMA_FAILED (8396L)
value ERROR_DS_REFERRAL (8235L)
value ERROR_DS_REFERRAL_LIMIT_EXCEEDED (8260L)
value ERROR_DS_REFUSING_FSMO_ROLES (8433L)
value ERROR_DS_REMOTE_CROSSREF_OP_FAILED (8601L)
value ERROR_DS_REPLICATOR_ONLY (8370L)
value ERROR_DS_REPLICA_SET_CHANGE_NOT_ALLOWED_ON_DISABLED_CR (8595L)
value ERROR_DS_REPL_LIFETIME_EXCEEDED (8614L)
value ERROR_DS_RESERVED_LINK_ID (8576L)
value ERROR_DS_RESERVED_MAPI_ID (8631L)
value ERROR_DS_RIDMGR_DISABLED (8263L)
value ERROR_DS_RIDMGR_INIT_ERROR (8211L)
value ERROR_DS_ROLE_NOT_VERIFIED (8610L)
value ERROR_DS_ROOT_CANT_BE_SUBREF (8326L)
value ERROR_DS_ROOT_MUST_BE_NC (8301L)
value ERROR_DS_ROOT_REQUIRES_CLASS_TOP (8432L)
value ERROR_DS_SAM_INIT_FAILURE (8504L)
value ERROR_DS_SAM_INIT_FAILURE_CONSOLE (8562L)
value ERROR_DS_SAM_NEED_BOOTKEY_FLOPPY (8530L)
value ERROR_DS_SAM_NEED_BOOTKEY_PASSWORD (8529L)
value ERROR_DS_SCHEMA_ALLOC_FAILED (8415L)
value ERROR_DS_SCHEMA_NOT_LOADED (8414L)
value ERROR_DS_SCHEMA_UPDATE_DISALLOWED (8509L)
value ERROR_DS_SECURITY_CHECKING_ERROR (8413L)
value ERROR_DS_SECURITY_ILLEGAL_MODIFY (8423L)
value ERROR_DS_SEC_DESC_INVALID (8354L)
value ERROR_DS_SEC_DESC_TOO_SHORT (8353L)
value ERROR_DS_SEMANTIC_ATT_TEST (8383L)
value ERROR_DS_SENSITIVE_GROUP_VIOLATION (8505L)
value ERROR_DS_SERVER_DOWN (8250L)
value ERROR_DS_SHUTTING_DOWN (8364L)
value ERROR_DS_SINGLE_USER_MODE_FAILED (8590L)
value ERROR_DS_SINGLE_VALUE_CONSTRAINT (8321L)
value ERROR_DS_SIZELIMIT_EXCEEDED (8227L)
value ERROR_DS_SORT_CONTROL_MISSING (8261L)
value ERROR_DS_SOURCE_AUDITING_NOT_ENABLED (8552L)
value ERROR_DS_SOURCE_DOMAIN_IN_FOREST (8534L)
value ERROR_DS_SPN_VALUE_NOT_UNIQUE_IN_FOREST (8647L)
value ERROR_DS_SRC_AND_DST_NC_IDENTICAL (8485L)
value ERROR_DS_SRC_AND_DST_OBJECT_CLASS_MISMATCH (8540L)
value ERROR_DS_SRC_GUID_MISMATCH (8488L)
value ERROR_DS_SRC_NAME_MISMATCH (8484L)
value ERROR_DS_SRC_OBJ_NOT_GROUP_OR_USER (8538L)
value ERROR_DS_SRC_SID_EXISTS_IN_FOREST (8539L)
value ERROR_DS_STRING_SD_CONVERSION_FAILED (8522L)
value ERROR_DS_STRONG_AUTH_REQUIRED (8232L)
value ERROR_DS_SUBREF_MUST_HAVE_PARENT (8356L)
value ERROR_DS_SUBTREE_NOTIFY_NOT_NC_HEAD (8376L)
value ERROR_DS_SUB_CLS_TEST_FAIL (8391L)
value ERROR_DS_SYNTAX_MISMATCH (8384L)
value ERROR_DS_THREAD_LIMIT_EXCEEDED (8587L)
value ERROR_DS_TIMELIMIT_EXCEEDED (8226L)
value ERROR_DS_TREE_DELETE_NOT_FINISHED (8397L)
value ERROR_DS_UNABLE_TO_SURRENDER_ROLES (8435L)
value ERROR_DS_UNAVAILABLE (8207L)
value ERROR_DS_UNAVAILABLE_CRIT_EXTENSION (8236L)
value ERROR_DS_UNDELETE_SAM_VALIDATION_FAILED (8645L)
value ERROR_DS_UNICODEPWD_NOT_IN_QUOTES (8556L)
value ERROR_DS_UNIVERSAL_CANT_HAVE_LOCAL_MEMBER (8518L)
value ERROR_DS_UNKNOWN_ERROR (8431L)
value ERROR_DS_UNKNOWN_OPERATION (8365L)
value ERROR_DS_UNWILLING_TO_PERFORM (8245L)
value ERROR_DS_UPN_VALUE_NOT_UNIQUE_IN_FOREST (8648L)
value ERROR_DS_USER_BUFFER_TO_SMALL (8309L)
value ERROR_DS_VALUE_KEY_NOT_UNIQUE (8650L)
value ERROR_DS_VERSION_CHECK_FAILURE (643L)
value ERROR_DS_WKO_CONTAINER_CANNOT_BE_SPECIAL (8611L)
value ERROR_DS_WRONG_LINKED_ATT_SYNTAX (8528L)
value ERROR_DS_WRONG_OM_OBJ_CLASS (8476L)
value ERROR_DUPLICATE_PRIVILEGES (311L)
value ERROR_DUPLICATE_SERVICE_NAME (1078L)
value ERROR_DUPLICATE_TAG (2014L)
value ERROR_DUP_DOMAINNAME (1221L)
value ERROR_DUP_NAME (52L)
value ERROR_DYNAMIC_CODE_BLOCKED (1655L)
value ERROR_DYNLINK_FROM_INVALID_RING (196L)
value ERROR_EAS_DIDNT_FIT (275L)
value ERROR_EAS_NOT_SUPPORTED (282L)
value ERROR_EA_ACCESS_DENIED (994L)
value ERROR_EA_FILE_CORRUPT (276L)
value ERROR_EA_LIST_INCONSISTENT (255L)
value ERROR_EA_TABLE_FULL (277L)
value ERROR_EC_CIRCULAR_FORWARDING (15082L)
value ERROR_EC_CREDSTORE_FULL (15083L)
value ERROR_EC_CRED_NOT_FOUND (15084L)
value ERROR_EC_LOG_DISABLED (15081L)
value ERROR_EC_NO_ACTIVE_CHANNEL (15085L)
value ERROR_EC_SUBSCRIPTION_CANNOT_ACTIVATE (15080L)
value ERROR_EDP_DPL_POLICY_CANT_BE_SATISFIED (357L)
value ERROR_EDP_POLICY_DENIES_OPERATION (356L)
value ERROR_EFS_ALG_BLOB_TOO_BIG (6013L)
value ERROR_EFS_DISABLED (6015L)
value ERROR_EFS_NOT_ALLOWED_IN_TRANSACTION (6831L)
value ERROR_EFS_SERVER_NOT_TRUSTED (6011L)
value ERROR_EFS_VERSION_NOT_SUPPORT (6016L)
value ERROR_ELEVATION_REQUIRED (740L)
value ERROR_EMPTY (4306L)
value ERROR_ENCLAVE_FAILURE (349L)
value ERROR_ENCLAVE_NOT_TERMINATED (814L)
value ERROR_ENCLAVE_VIOLATION (815L)
value ERROR_ENCRYPTED_FILE_NOT_SUPPORTED (489L)
value ERROR_ENCRYPTED_IO_NOT_POSSIBLE (808L)
value ERROR_ENCRYPTING_METADATA_DISALLOWED (431L)
value ERROR_ENCRYPTION_DISABLED (430L)
value ERROR_ENCRYPTION_FAILED (6000L)
value ERROR_ENCRYPTION_POLICY_DENIES_OPERATION (6022L)
value ERROR_END_OF_MEDIA (1100L)
value ERROR_ENLISTMENT_NOT_FOUND (6717L)
value ERROR_ENLISTMENT_NOT_SUPERIOR (6820L)
value ERROR_ENVVAR_NOT_FOUND (203L)
value ERROR_EOM_OVERFLOW (1129L)
value ERROR_ERRORS_ENCOUNTERED (774L)
value ERROR_EVALUATION_EXPIRATION (622L)
value ERROR_EVENTLOG_CANT_START (1501L)
value ERROR_EVENTLOG_FILE_CHANGED (1503L)
value ERROR_EVENTLOG_FILE_CORRUPT (1500L)
value ERROR_EVENT_DONE (710L)
value ERROR_EVENT_PENDING (711L)
value ERROR_EVT_CANNOT_OPEN_CHANNEL_OF_QUERY (15036L)
value ERROR_EVT_CHANNEL_CANNOT_ACTIVATE (15025L)
value ERROR_EVT_CHANNEL_NOT_FOUND (15007L)
value ERROR_EVT_CONFIGURATION_ERROR (15010L)
value ERROR_EVT_EVENT_DEFINITION_NOT_FOUND (15032L)
value ERROR_EVT_EVENT_TEMPLATE_NOT_FOUND (15003L)
value ERROR_EVT_FILTER_ALREADYSCOPED (15014L)
value ERROR_EVT_FILTER_INVARG (15016L)
value ERROR_EVT_FILTER_INVTEST (15017L)
value ERROR_EVT_FILTER_INVTYPE (15018L)
value ERROR_EVT_FILTER_NOTELTSET (15015L)
value ERROR_EVT_FILTER_OUT_OF_RANGE (15038L)
value ERROR_EVT_FILTER_PARSEERR (15019L)
value ERROR_EVT_FILTER_TOO_COMPLEX (15026L)
value ERROR_EVT_FILTER_UNEXPECTEDTOKEN (15021L)
value ERROR_EVT_FILTER_UNSUPPORTEDOP (15020L)
value ERROR_EVT_INVALID_CHANNEL_PATH (15000L)
value ERROR_EVT_INVALID_CHANNEL_PROPERTY_VALUE (15023L)
value ERROR_EVT_INVALID_EVENT_DATA (15005L)
value ERROR_EVT_INVALID_OPERATION_OVER_ENABLED_DIRECT_CHANNEL (15022L)
value ERROR_EVT_INVALID_PUBLISHER_NAME (15004L)
value ERROR_EVT_INVALID_PUBLISHER_PROPERTY_VALUE (15024L)
value ERROR_EVT_INVALID_QUERY (15001L)
value ERROR_EVT_MALFORMED_XML_TEXT (15008L)
value ERROR_EVT_MAX_INSERTS_REACHED (15031L)
value ERROR_EVT_MESSAGE_ID_NOT_FOUND (15028L)
value ERROR_EVT_MESSAGE_LOCALE_NOT_FOUND (15033L)
value ERROR_EVT_MESSAGE_NOT_FOUND (15027L)
value ERROR_EVT_NON_VALIDATING_MSXML (15013L)
value ERROR_EVT_PUBLISHER_DISABLED (15037L)
value ERROR_EVT_PUBLISHER_METADATA_NOT_FOUND (15002L)
value ERROR_EVT_QUERY_RESULT_INVALID_POSITION (15012L)
value ERROR_EVT_QUERY_RESULT_STALE (15011L)
value ERROR_EVT_SUBSCRIPTION_TO_DIRECT_CHANNEL (15009L)
value ERROR_EVT_UNRESOLVED_PARAMETER_INSERT (15030L)
value ERROR_EVT_UNRESOLVED_VALUE_INSERT (15029L)
value ERROR_EVT_VERSION_TOO_NEW (15035L)
value ERROR_EVT_VERSION_TOO_OLD (15034L)
value ERROR_EXCEPTION_IN_RESOURCE_CALL (5930L)
value ERROR_EXCEPTION_IN_SERVICE (1064L)
value ERROR_EXCL_SEM_ALREADY_OWNED (101L)
value ERROR_EXE_CANNOT_MODIFY_SIGNED_BINARY (217L)
value ERROR_EXE_CANNOT_MODIFY_STRONG_SIGNED_BINARY (218L)
value ERROR_EXE_MACHINE_TYPE_MISMATCH (216L)
value ERROR_EXE_MARKED_INVALID (192L)
value ERROR_EXPIRED_HANDLE (6854L)
value ERROR_EXTENDED_ERROR (1208L)
value ERROR_EXTERNAL_BACKING_PROVIDER_UNKNOWN (343L)
value ERROR_EXTERNAL_SYSKEY_NOT_SUPPORTED (399L)
value ERROR_EXTRANEOUS_INFORMATION (677L)
value ERROR_FAILED_DRIVER_ENTRY (647L)
value ERROR_FAILED_SERVICE_CONTROLLER_CONNECT (1063L)
value ERROR_FAIL_FAST_EXCEPTION (1653L)
value ERROR_FAIL_NOACTION_REBOOT (350L)
value ERROR_FAIL_REBOOT_INITIATED (3018L)
value ERROR_FAIL_REBOOT_REQUIRED (3017L)
value ERROR_FAIL_RESTART (352L)
value ERROR_FAIL_SHUTDOWN (351L)
value ERROR_FATAL_APP_EXIT (713L)
value ERROR_FILEMARK_DETECTED (1101L)
value ERROR_FILENAME_EXCED_RANGE (206L)
value ERROR_FILE_CHECKED_OUT (220L)
value ERROR_FILE_CORRUPT (1392L)
value ERROR_FILE_ENCRYPTED (6002L)
value ERROR_FILE_EXISTS (80L)
value ERROR_FILE_HANDLE_REVOKED (806L)
value ERROR_FILE_IDENTITY_NOT_PERSISTENT (6823L)
value ERROR_FILE_INVALID (1006L)
value ERROR_FILE_LEVEL_TRIM_NOT_SUPPORTED (326L)
value ERROR_FILE_METADATA_OPTIMIZATION_IN_PROGRESS (809L)
value ERROR_FILE_NOT_ENCRYPTED (6007L)
value ERROR_FILE_NOT_FOUND (2L)
value ERROR_FILE_NOT_SUPPORTED (425L)
value ERROR_FILE_OFFLINE (4350L)
value ERROR_FILE_PROTECTED_UNDER_DPL (406L)
value ERROR_FILE_READ_ONLY (6009L)
value ERROR_FILE_SHARE_RESOURCE_CONFLICT (5938L)
value ERROR_FILE_SNAP_INVALID_PARAMETER (440L)
value ERROR_FILE_SNAP_IN_PROGRESS (435L)
value ERROR_FILE_SNAP_IO_NOT_COORDINATED (438L)
value ERROR_FILE_SNAP_MODIFY_NOT_SUPPORTED (437L)
value ERROR_FILE_SNAP_UNEXPECTED_ERROR (439L)
value ERROR_FILE_SNAP_USER_SECTION_NOT_SUPPORTED (436L)
value ERROR_FILE_SYSTEM_LIMITATION (665L)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_BUSY (371L)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_INVALID_OPERATION (385L)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_METADATA_CORRUPT (370L)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_PROVIDER_UNKNOWN (372L)
value ERROR_FILE_SYSTEM_VIRTUALIZATION_UNAVAILABLE (369L)
value ERROR_FILE_TOO_LARGE (223L)
value ERROR_FIRMWARE_UPDATED (728L)
value ERROR_FLOATED_SECTION (6846L)
value ERROR_FLOAT_MULTIPLE_FAULTS (630L)
value ERROR_FLOAT_MULTIPLE_TRAPS (631L)
value ERROR_FLOPPY_BAD_REGISTERS (1125L)
value ERROR_FLOPPY_ID_MARK_NOT_FOUND (1122L)
value ERROR_FLOPPY_UNKNOWN_ERROR (1124L)
value ERROR_FLOPPY_VOLUME (584L)
value ERROR_FLOPPY_WRONG_CYLINDER (1123L)
value ERROR_FORMS_AUTH_REQUIRED (224L)
value ERROR_FOUND_OUT_OF_SCOPE (601L)
value ERROR_FSFILTER_OP_COMPLETED_SUCCESSFULLY (762L)
value ERROR_FS_DRIVER_REQUIRED (588L)
value ERROR_FS_METADATA_INCONSISTENT (510L)
value ERROR_FT_DI_SCAN_REQUIRED (339L)
value ERROR_FT_READ_FAILURE (415L)
value ERROR_FT_READ_FROM_COPY_FAILURE (818L)
value ERROR_FT_READ_RECOVERY_FROM_BACKUP (704L)
value ERROR_FT_WRITE_FAILURE (338L)
value ERROR_FT_WRITE_RECOVERY (705L)
value ERROR_FULLSCREEN_MODE (1007L)
value ERROR_FULL_BACKUP (4004L)
value ERROR_FUNCTION_FAILED (1627L)
value ERROR_FUNCTION_NOT_CALLED (1626L)
value ERROR_GDI_HANDLE_LEAK (373L)
value ERROR_GENERIC_COMMAND_FAILED (14109L)
value ERROR_GENERIC_NOT_MAPPED (1360L)
value ERROR_GEN_FAILURE (31L)
value ERROR_GLOBAL_ONLY_HOOK (1429L)
value ERROR_GPIO_CLIENT_INFORMATION_INVALID (15322L)
value ERROR_GPIO_INCOMPATIBLE_CONNECT_MODE (15326L)
value ERROR_GPIO_INTERRUPT_ALREADY_UNMASKED (15327L)
value ERROR_GPIO_INVALID_REGISTRATION_PACKET (15324L)
value ERROR_GPIO_OPERATION_DENIED (15325L)
value ERROR_GPIO_VERSION_NOT_SUPPORTED (15323L)
value ERROR_GRACEFUL_DISCONNECT (1226L)
value ERROR_GROUPSET_CANT_PROVIDE (5993L)
value ERROR_GROUPSET_NOT_AVAILABLE (5991L)
value ERROR_GROUPSET_NOT_FOUND (5992L)
value ERROR_GROUP_EXISTS (1318L)
value ERROR_GROUP_NOT_AVAILABLE (5012L)
value ERROR_GROUP_NOT_FOUND (5013L)
value ERROR_GROUP_NOT_ONLINE (5014L)
value ERROR_GUID_SUBSTITUTION_MADE (680L)
value ERROR_HANDLES_CLOSED (676L)
value ERROR_HANDLE_DISK_FULL (39L)
value ERROR_HANDLE_EOF (38L)
value ERROR_HANDLE_NO_LONGER_VALID (6815L)
value ERROR_HANDLE_REVOKED (811L)
value ERROR_HASH_NOT_PRESENT (15301L)
value ERROR_HASH_NOT_SUPPORTED (15300L)
value ERROR_HAS_SYSTEM_CRITICAL_FILES (488L)
value ERROR_HEURISTIC_DAMAGE_POSSIBLE (6731L)
value ERROR_HIBERNATED (726L)
value ERROR_HIBERNATION_FAILURE (656L)
value ERROR_HISTORY_DIRECTORY_ENTRY_DEFAULT_COUNT (8)
value ERROR_HOOK_NEEDS_HMOD (1428L)
value ERROR_HOOK_NOT_INSTALLED (1431L)
value ERROR_HOOK_TYPE_NOT_ALLOWED (1458L)
value ERROR_HOST_DOWN (1256L)
value ERROR_HOST_NODE_NOT_AVAILABLE (5005L)
value ERROR_HOST_NODE_NOT_GROUP_OWNER (5016L)
value ERROR_HOST_NODE_NOT_RESOURCE_OWNER (5015L)
value ERROR_HOST_UNREACHABLE (1232L)
value ERROR_HOTKEY_ALREADY_REGISTERED (1409L)
value ERROR_HOTKEY_NOT_REGISTERED (1419L)
value ERROR_HWNDS_HAVE_DIFF_PARENT (1441L)
value ERROR_ICM_NOT_ENABLED (2018L)
value ERROR_IEPORT_FULL (4341L)
value ERROR_ILLEGAL_CHARACTER (582L)
value ERROR_ILLEGAL_DLL_RELOCATION (623L)
value ERROR_ILLEGAL_ELEMENT_ADDRESS (1162L)
value ERROR_ILLEGAL_FLOAT_CONTEXT (579L)
value ERROR_ILL_FORMED_PASSWORD (1324L)
value ERROR_IMAGE_AT_DIFFERENT_BASE (807L)
value ERROR_IMAGE_MACHINE_TYPE_MISMATCH (706L)
value ERROR_IMAGE_MACHINE_TYPE_MISMATCH_EXE (720L)
value ERROR_IMAGE_NOT_AT_BASE (700L)
value ERROR_IMAGE_SUBSYSTEM_NOT_PRESENT (308L)
value ERROR_IMPLEMENTATION_LIMIT (1292L)
value ERROR_IMPLICIT_TRANSACTION_NOT_SUPPORTED (6725L)
value ERROR_INCOMPATIBLE_SERVICE_PRIVILEGE (1297L)
value ERROR_INCOMPATIBLE_SERVICE_SID_TYPE (1290L)
value ERROR_INCOMPATIBLE_WITH_GLOBAL_SHORT_NAME_REGISTRY_SETTING (304L)
value ERROR_INCORRECT_ACCOUNT_TYPE (8646L)
value ERROR_INCORRECT_ADDRESS (1241L)
value ERROR_INCORRECT_SIZE (1462L)
value ERROR_INC_BACKUP (4003L)
value ERROR_INDEX_ABSENT (1611L)
value ERROR_INDEX_OUT_OF_BOUNDS (474L)
value ERROR_INDIGENOUS_TYPE (4338L)
value ERROR_INDOUBT_TRANSACTIONS_EXIST (6827L)
value ERROR_INFLOOP_IN_RELOC_CHAIN (202L)
value ERROR_INSTALL_ALREADY_RUNNING (1618L)
value ERROR_INSTALL_CANCEL (15608L)
value ERROR_INSTALL_DEREGISTRATION_FAILURE (15607L)
value ERROR_INSTALL_FAILED (15609L)
value ERROR_INSTALL_FAILURE (1603L)
value ERROR_INSTALL_FIREWALL_SERVICE_NOT_RUNNING (15626L)
value ERROR_INSTALL_FULLTRUST_HOSTRUNTIME_REQUIRES_MAIN_PACKAGE_FULLTRUST_CAPABILITY (15663L)
value ERROR_INSTALL_INVALID_PACKAGE (15602L)
value ERROR_INSTALL_INVALID_RELATED_SET_UPDATE (15639L)
value ERROR_INSTALL_LANGUAGE_UNSUPPORTED (1623L)
value ERROR_INSTALL_LOG_FAILURE (1622L)
value ERROR_INSTALL_NETWORK_FAILURE (15605L)
value ERROR_INSTALL_NOTUSED (1634L)
value ERROR_INSTALL_OPEN_PACKAGE_FAILED (15600L)
value ERROR_INSTALL_OPTIONAL_PACKAGE_APPLICATIONID_NOT_UNIQUE (15637L)
value ERROR_INSTALL_OPTIONAL_PACKAGE_REQUIRES_MAIN_PACKAGE (15634L)
value ERROR_INSTALL_OPTIONAL_PACKAGE_REQUIRES_MAIN_PACKAGE_FULLTRUST_CAPABILITY (15640L)
value ERROR_INSTALL_OUT_OF_DISK_SPACE (15604L)
value ERROR_INSTALL_PACKAGE_DOWNGRADE (15622L)
value ERROR_INSTALL_PACKAGE_INVALID (1620L)
value ERROR_INSTALL_PACKAGE_NOT_FOUND (15601L)
value ERROR_INSTALL_PACKAGE_OPEN_FAILED (1619L)
value ERROR_INSTALL_PACKAGE_REJECTED (1625L)
value ERROR_INSTALL_PACKAGE_VERSION (1613L)
value ERROR_INSTALL_PLATFORM_UNSUPPORTED (1633L)
value ERROR_INSTALL_POLICY_FAILURE (15615L)
value ERROR_INSTALL_PREREQUISITE_FAILED (15613L)
value ERROR_INSTALL_REGISTRATION_FAILURE (15606L)
value ERROR_INSTALL_REJECTED (1654L)
value ERROR_INSTALL_REMOTE_DISALLOWED (1640L)
value ERROR_INSTALL_REMOTE_PROHIBITED (1645L)
value ERROR_INSTALL_RESOLVE_DEPENDENCY_FAILED (15603L)
value ERROR_INSTALL_RESOLVE_HOSTRUNTIME_DEPENDENCY_FAILED (15665L)
value ERROR_INSTALL_SERVICE_FAILURE (1601L)
value ERROR_INSTALL_SERVICE_SAFEBOOT (1652L)
value ERROR_INSTALL_SOURCE_ABSENT (1612L)
value ERROR_INSTALL_SUSPEND (1604L)
value ERROR_INSTALL_TEMP_UNWRITABLE (1632L)
value ERROR_INSTALL_TRANSFORM_FAILURE (1624L)
value ERROR_INSTALL_TRANSFORM_REJECTED (1644L)
value ERROR_INSTALL_UI_FAILURE (1621L)
value ERROR_INSTALL_USEREXIT (1602L)
value ERROR_INSTALL_VOLUME_CORRUPT (15630L)
value ERROR_INSTALL_VOLUME_NOT_EMPTY (15628L)
value ERROR_INSTALL_VOLUME_OFFLINE (15629L)
value ERROR_INSTALL_WRONG_PROCESSOR_ARCHITECTURE (15632L)
value ERROR_INSTRUCTION_MISALIGNMENT (549L)
value ERROR_INSUFFICIENT_BUFFER (122L)
value ERROR_INSUFFICIENT_LOGON_INFO (608L)
value ERROR_INSUFFICIENT_POWER (639L)
value ERROR_INSUFFICIENT_RESOURCE_FOR_SPECIFIED_SHARED_SECTION_SIZE (781L)
value ERROR_INSUFFICIENT_VIRTUAL_ADDR_RESOURCES (473L)
value ERROR_INTERMIXED_KERNEL_EA_OPERATION (324L)
value ERROR_INTERNAL_DB_CORRUPTION (1358L)
value ERROR_INTERNAL_DB_ERROR (1383L)
value ERROR_INTERNAL_ERROR (1359L)
value ERROR_INTERRUPT_STILL_CONNECTED (764L)
value ERROR_INTERRUPT_VECTOR_ALREADY_CONNECTED (763L)
value ERROR_INVALID_ACCEL_HANDLE (1403L)
value ERROR_INVALID_ACCESS (12L)
value ERROR_INVALID_ACCOUNT_NAME (1315L)
value ERROR_INVALID_ACE_CONDITION (805L)
value ERROR_INVALID_ACL (1336L)
value ERROR_INVALID_ADDRESS (487L)
value ERROR_INVALID_AT_INTERRUPT_TIME (104L)
value ERROR_INVALID_BLOCK (9L)
value ERROR_INVALID_BLOCK_LENGTH (1106L)
value ERROR_INVALID_CAP (320L)
value ERROR_INVALID_CATEGORY (117L)
value ERROR_INVALID_CLEANER (4310L)
value ERROR_INVALID_CMM (2010L)
value ERROR_INVALID_COLORINDEX (2022L)
value ERROR_INVALID_COLORSPACE (2017L)
value ERROR_INVALID_COMBOBOX_MESSAGE (1422L)
value ERROR_INVALID_COMMAND_LINE (1639L)
value ERROR_INVALID_COMPUTERNAME (1210L)
value ERROR_INVALID_CRUNTIME_PARAMETER (1288L)
value ERROR_INVALID_CURSOR_HANDLE (1402L)
value ERROR_INVALID_DATA (13L)
value ERROR_INVALID_DATATYPE (1804L)
value ERROR_INVALID_DEVICE_OBJECT_PARAMETER (650L)
value ERROR_INVALID_DLL (1154L)
value ERROR_INVALID_DOMAINNAME (1212L)
value ERROR_INVALID_DOMAIN_ROLE (1354L)
value ERROR_INVALID_DOMAIN_STATE (1353L)
value ERROR_INVALID_DRIVE (15L)
value ERROR_INVALID_DRIVE_OBJECT (4321L)
value ERROR_INVALID_DWP_HANDLE (1405L)
value ERROR_INVALID_EA_HANDLE (278L)
value ERROR_INVALID_EA_NAME (254L)
value ERROR_INVALID_EDIT_HEIGHT (1424L)
value ERROR_INVALID_ENVIRONMENT (1805L)
value ERROR_INVALID_EVENTNAME (1211L)
value ERROR_INVALID_EVENT_COUNT (151L)
value ERROR_INVALID_EXCEPTION_HANDLER (310L)
value ERROR_INVALID_EXE_SIGNATURE (191L)
value ERROR_INVALID_FIELD (1616L)
value ERROR_INVALID_FIELD_IN_PARAMETER_LIST (328L)
value ERROR_INVALID_FILTER_PROC (1427L)
value ERROR_INVALID_FLAGS (1004L)
value ERROR_INVALID_FLAG_NUMBER (186L)
value ERROR_INVALID_FORM_NAME (1902L)
value ERROR_INVALID_FORM_SIZE (1903L)
value ERROR_INVALID_FUNCTION (1L)
value ERROR_INVALID_GROUPNAME (1209L)
value ERROR_INVALID_GROUP_ATTRIBUTES (1345L)
value ERROR_INVALID_GW_COMMAND (1443L)
value ERROR_INVALID_HANDLE (6L)
value ERROR_INVALID_HANDLE_STATE (1609L)
value ERROR_INVALID_HOOK_FILTER (1426L)
value ERROR_INVALID_HOOK_HANDLE (1404L)
value ERROR_INVALID_HW_PROFILE (619L)
value ERROR_INVALID_ICON_HANDLE (1414L)
value ERROR_INVALID_ID_AUTHORITY (1343L)
value ERROR_INVALID_IMAGE_HASH (577L)
value ERROR_INVALID_IMPORT_OF_NON_DLL (1276L)
value ERROR_INVALID_INDEX (1413L)
value ERROR_INVALID_KERNEL_INFO_VERSION (340L)
value ERROR_INVALID_KEYBOARD_HANDLE (1457L)
value ERROR_INVALID_LABEL (1299L)
value ERROR_INVALID_LB_MESSAGE (1432L)
value ERROR_INVALID_LDT_DESCRIPTOR (564L)
value ERROR_INVALID_LDT_OFFSET (563L)
value ERROR_INVALID_LDT_SIZE (561L)
value ERROR_INVALID_LEVEL (124L)
value ERROR_INVALID_LIBRARY (4301L)
value ERROR_INVALID_LIST_FORMAT (153L)
value ERROR_INVALID_LOCK_RANGE (307L)
value ERROR_INVALID_LOGON_HOURS (1328L)
value ERROR_INVALID_LOGON_TYPE (1367L)
value ERROR_INVALID_MEDIA (4300L)
value ERROR_INVALID_MEDIA_POOL (4302L)
value ERROR_INVALID_MEMBER (1388L)
value ERROR_INVALID_MENU_HANDLE (1401L)
value ERROR_INVALID_MESSAGE (1002L)
value ERROR_INVALID_MESSAGEDEST (1218L)
value ERROR_INVALID_MESSAGENAME (1217L)
value ERROR_INVALID_MINALLOCSIZE (195L)
value ERROR_INVALID_MODULETYPE (190L)
value ERROR_INVALID_MONITOR_HANDLE (1461L)
value ERROR_INVALID_MSGBOX_STYLE (1438L)
value ERROR_INVALID_NAME (123L)
value ERROR_INVALID_NETNAME (1214L)
value ERROR_INVALID_OPERATION (4317L)
value ERROR_INVALID_OPERATION_ON_QUORUM (5068L)
value ERROR_INVALID_OPLOCK_PROTOCOL (301L)
value ERROR_INVALID_ORDINAL (182L)
value ERROR_INVALID_OWNER (1307L)
value ERROR_INVALID_PACKAGE_SID_LENGTH (4253L)
value ERROR_INVALID_PARAMETER (87L)
value ERROR_INVALID_PASSWORD (86L)
value ERROR_INVALID_PASSWORDNAME (1216L)
value ERROR_INVALID_PATCH_XML (1650L)
value ERROR_INVALID_PEP_INFO_VERSION (341L)
value ERROR_INVALID_PIXEL_FORMAT (2000L)
value ERROR_INVALID_PLUGPLAY_DEVICE_PATH (620L)
value ERROR_INVALID_PORT_ATTRIBUTES (545L)
value ERROR_INVALID_PRIMARY_GROUP (1308L)
value ERROR_INVALID_PRINTER_COMMAND (1803L)
value ERROR_INVALID_PRINTER_DRIVER_MANIFEST (3021L)
value ERROR_INVALID_PRINTER_NAME (1801L)
value ERROR_INVALID_PRINTER_STATE (1906L)
value ERROR_INVALID_PRINT_MONITOR (3007L)
value ERROR_INVALID_PRIORITY (1800L)
value ERROR_INVALID_PROFILE (2011L)
value ERROR_INVALID_QUOTA_LOWER (547L)
value ERROR_INVALID_REPARSE_DATA (4392L)
value ERROR_INVALID_RUNLEVEL_SETTING (15401L)
value ERROR_INVALID_SCROLLBAR_RANGE (1448L)
value ERROR_INVALID_SECURITY_DESCR (1338L)
value ERROR_INVALID_SEGDPL (198L)
value ERROR_INVALID_SEGMENT_NUMBER (180L)
value ERROR_INVALID_SEPARATOR_FILE (1799L)
value ERROR_INVALID_SERVER_STATE (1352L)
value ERROR_INVALID_SERVICENAME (1213L)
value ERROR_INVALID_SERVICE_ACCOUNT (1057L)
value ERROR_INVALID_SERVICE_CONTROL (1052L)
value ERROR_INVALID_SERVICE_LOCK (1071L)
value ERROR_INVALID_SHARENAME (1215L)
value ERROR_INVALID_SHOWWIN_COMMAND (1449L)
value ERROR_INVALID_SID (1337L)
value ERROR_INVALID_SIGNAL_NUMBER (209L)
value ERROR_INVALID_SPI_VALUE (1439L)
value ERROR_INVALID_STACKSEG (189L)
value ERROR_INVALID_STAGED_SIGNATURE (15620L)
value ERROR_INVALID_STARTING_CODESEG (188L)
value ERROR_INVALID_STATE (5023L)
value ERROR_INVALID_SUB_AUTHORITY (1335L)
value ERROR_INVALID_TABLE (1628L)
value ERROR_INVALID_TARGET_HANDLE (114L)
value ERROR_INVALID_TASK_INDEX (1551L)
value ERROR_INVALID_TASK_NAME (1550L)
value ERROR_INVALID_THREAD_ID (1444L)
value ERROR_INVALID_TIME (1901L)
value ERROR_INVALID_TOKEN (315L)
value ERROR_INVALID_TRANSACTION (6700L)
value ERROR_INVALID_TRANSFORM (2020L)
value ERROR_INVALID_UNWIND_TARGET (544L)
value ERROR_INVALID_USER_BUFFER (1784L)
value ERROR_INVALID_USER_PRINCIPAL_NAME (8636L)
value ERROR_INVALID_VARIANT (604L)
value ERROR_INVALID_VERIFY_SWITCH (118L)
value ERROR_INVALID_WINDOW_HANDLE (1400L)
value ERROR_INVALID_WINDOW_STYLE (2002L)
value ERROR_INVALID_WORKSTATION (1329L)
value ERROR_IOPL_NOT_ENABLED (197L)
value ERROR_IO_DEVICE (1117L)
value ERROR_IO_INCOMPLETE (996L)
value ERROR_IO_PENDING (997L)
value ERROR_IO_PRIVILEGE_FAILED (571L)
value ERROR_IO_REISSUE_AS_CACHED (3950L)
value ERROR_IPSEC_AUTH_FIREWALL_DROP (13917L)
value ERROR_IPSEC_BAD_SPI (13910L)
value ERROR_IPSEC_CLEAR_TEXT_DROP (13916L)
value ERROR_IPSEC_DEFAULT_MM_AUTH_NOT_FOUND (13014L)
value ERROR_IPSEC_DEFAULT_MM_POLICY_NOT_FOUND (13013L)
value ERROR_IPSEC_DEFAULT_QM_POLICY_NOT_FOUND (13015L)
value ERROR_IPSEC_DOSP_BLOCK (13925L)
value ERROR_IPSEC_DOSP_INVALID_PACKET (13927L)
value ERROR_IPSEC_DOSP_KEYMOD_NOT_ALLOWED (13930L)
value ERROR_IPSEC_DOSP_MAX_ENTRIES (13929L)
value ERROR_IPSEC_DOSP_MAX_PER_IP_RATELIMIT_QUEUES (13932L)
value ERROR_IPSEC_DOSP_NOT_INSTALLED (13931L)
value ERROR_IPSEC_DOSP_RECEIVED_MULTICAST (13926L)
value ERROR_IPSEC_DOSP_STATE_LOOKUP_FAILED (13928L)
value ERROR_IPSEC_IKE_ADD_UPDATE_KEY_FAILED (13860L)
value ERROR_IPSEC_IKE_ATTRIB_FAIL (13802L)
value ERROR_IPSEC_IKE_AUTHORIZATION_FAILURE (13905L)
value ERROR_IPSEC_IKE_AUTHORIZATION_FAILURE_WITH_OPTIONAL_RETRY (13907L)
value ERROR_IPSEC_IKE_AUTH_FAIL (13801L)
value ERROR_IPSEC_IKE_BENIGN_REINIT (13878L)
value ERROR_IPSEC_IKE_CERT_CHAIN_POLICY_MISMATCH (13887L)
value ERROR_IPSEC_IKE_CGA_AUTH_FAILED (13892L)
value ERROR_IPSEC_IKE_COEXISTENCE_SUPPRESS (13902L)
value ERROR_IPSEC_IKE_CRITICAL_PAYLOAD_NOT_RECOGNIZED (13823L)
value ERROR_IPSEC_IKE_CRL_FAILED (13817L)
value ERROR_IPSEC_IKE_DECRYPT (13867L)
value ERROR_IPSEC_IKE_DH_FAIL (13822L)
value ERROR_IPSEC_IKE_DH_FAILURE (13864L)
value ERROR_IPSEC_IKE_DOS_COOKIE_SENT (13890L)
value ERROR_IPSEC_IKE_DROP_NO_RESPONSE (13813L)
value ERROR_IPSEC_IKE_ENCRYPT (13866L)
value ERROR_IPSEC_IKE_ERROR (13816L)
value ERROR_IPSEC_IKE_FAILQUERYSSP (13854L)
value ERROR_IPSEC_IKE_FAILSSPINIT (13853L)
value ERROR_IPSEC_IKE_GENERAL_PROCESSING_ERROR (13804L)
value ERROR_IPSEC_IKE_GETSPIFAIL (13857L)
value ERROR_IPSEC_IKE_INNER_IP_ASSIGNMENT_FAILURE (13899L)
value ERROR_IPSEC_IKE_INVALID_AUTH_ALG (13874L)
value ERROR_IPSEC_IKE_INVALID_AUTH_PAYLOAD (13889L)
value ERROR_IPSEC_IKE_INVALID_CERT_KEYLEN (13881L)
value ERROR_IPSEC_IKE_INVALID_CERT_TYPE (13819L)
value ERROR_IPSEC_IKE_INVALID_COOKIE (13846L)
value ERROR_IPSEC_IKE_INVALID_ENCRYPT_ALG (13873L)
value ERROR_IPSEC_IKE_INVALID_FILTER (13858L)
value ERROR_IPSEC_IKE_INVALID_GROUP (13865L)
value ERROR_IPSEC_IKE_INVALID_HASH (13870L)
value ERROR_IPSEC_IKE_INVALID_HASH_ALG (13871L)
value ERROR_IPSEC_IKE_INVALID_HASH_SIZE (13872L)
value ERROR_IPSEC_IKE_INVALID_HEADER (13824L)
value ERROR_IPSEC_IKE_INVALID_KEY_USAGE (13818L)
value ERROR_IPSEC_IKE_INVALID_MAJOR_VERSION (13880L)
value ERROR_IPSEC_IKE_INVALID_MM_FOR_QM (13894L)
value ERROR_IPSEC_IKE_INVALID_PAYLOAD (13843L)
value ERROR_IPSEC_IKE_INVALID_POLICY (13861L)
value ERROR_IPSEC_IKE_INVALID_RESPONDER_LIFETIME_NOTIFY (13879L)
value ERROR_IPSEC_IKE_INVALID_SIG (13875L)
value ERROR_IPSEC_IKE_INVALID_SIGNATURE (13826L)
value ERROR_IPSEC_IKE_INVALID_SITUATION (13863L)
value ERROR_IPSEC_IKE_KERBEROS_ERROR (13827L)
value ERROR_IPSEC_IKE_KILL_DUMMY_NAP_TUNNEL (13898L)
value ERROR_IPSEC_IKE_LOAD_FAILED (13876L)
value ERROR_IPSEC_IKE_LOAD_SOFT_SA (13844L)
value ERROR_IPSEC_IKE_MM_ACQUIRE_DROP (13809L)
value ERROR_IPSEC_IKE_MM_DELAY_DROP (13814L)
value ERROR_IPSEC_IKE_MM_EXPIRED (13885L)
value ERROR_IPSEC_IKE_MM_LIMIT (13882L)
value ERROR_IPSEC_IKE_NEGOTIATION_DISABLED (13883L)
value ERROR_IPSEC_IKE_NEGOTIATION_PENDING (13803L)
value ERROR_IPSEC_IKE_NEG_STATUS_BEGIN (13800L)
value ERROR_IPSEC_IKE_NEG_STATUS_END (13897L)
value ERROR_IPSEC_IKE_NEG_STATUS_EXTENDED_END (13909L)
value ERROR_IPSEC_IKE_NOTCBPRIV (13851L)
value ERROR_IPSEC_IKE_NO_CERT (13806L)
value ERROR_IPSEC_IKE_NO_MM_POLICY (13850L)
value ERROR_IPSEC_IKE_NO_PEER_CERT (13847L)
value ERROR_IPSEC_IKE_NO_POLICY (13825L)
value ERROR_IPSEC_IKE_NO_PRIVATE_KEY (13820L)
value ERROR_IPSEC_IKE_NO_PUBLIC_KEY (13828L)
value ERROR_IPSEC_IKE_OUT_OF_MEMORY (13859L)
value ERROR_IPSEC_IKE_PEER_CRL_FAILED (13848L)
value ERROR_IPSEC_IKE_PEER_DOESNT_SUPPORT_MOBIKE (13904L)
value ERROR_IPSEC_IKE_PEER_MM_ASSUMED_INVALID (13886L)
value ERROR_IPSEC_IKE_POLICY_CHANGE (13849L)
value ERROR_IPSEC_IKE_POLICY_MATCH (13868L)
value ERROR_IPSEC_IKE_PROCESS_ERR (13829L)
value ERROR_IPSEC_IKE_PROCESS_ERR_CERT (13835L)
value ERROR_IPSEC_IKE_PROCESS_ERR_CERT_REQ (13836L)
value ERROR_IPSEC_IKE_PROCESS_ERR_DELETE (13841L)
value ERROR_IPSEC_IKE_PROCESS_ERR_HASH (13837L)
value ERROR_IPSEC_IKE_PROCESS_ERR_ID (13834L)
value ERROR_IPSEC_IKE_PROCESS_ERR_KE (13833L)
value ERROR_IPSEC_IKE_PROCESS_ERR_NATOA (13893L)
value ERROR_IPSEC_IKE_PROCESS_ERR_NONCE (13839L)
value ERROR_IPSEC_IKE_PROCESS_ERR_NOTIFY (13840L)
value ERROR_IPSEC_IKE_PROCESS_ERR_PROP (13831L)
value ERROR_IPSEC_IKE_PROCESS_ERR_SA (13830L)
value ERROR_IPSEC_IKE_PROCESS_ERR_SIG (13838L)
value ERROR_IPSEC_IKE_PROCESS_ERR_TRANS (13832L)
value ERROR_IPSEC_IKE_PROCESS_ERR_VENDOR (13842L)
value ERROR_IPSEC_IKE_QM_ACQUIRE_DROP (13810L)
value ERROR_IPSEC_IKE_QM_DELAY_DROP (13815L)
value ERROR_IPSEC_IKE_QM_EXPIRED (13895L)
value ERROR_IPSEC_IKE_QM_LIMIT (13884L)
value ERROR_IPSEC_IKE_QUEUE_DROP_MM (13811L)
value ERROR_IPSEC_IKE_QUEUE_DROP_NO_MM (13812L)
value ERROR_IPSEC_IKE_RATELIMIT_DROP (13903L)
value ERROR_IPSEC_IKE_REQUIRE_CP_PAYLOAD_MISSING (13900L)
value ERROR_IPSEC_IKE_RPC_DELETE (13877L)
value ERROR_IPSEC_IKE_SA_DELETED (13807L)
value ERROR_IPSEC_IKE_SA_REAPED (13808L)
value ERROR_IPSEC_IKE_SECLOADFAIL (13852L)
value ERROR_IPSEC_IKE_SHUTTING_DOWN (13891L)
value ERROR_IPSEC_IKE_SIMULTANEOUS_REKEY (13821L)
value ERROR_IPSEC_IKE_SOFT_SA_TORN_DOWN (13845L)
value ERROR_IPSEC_IKE_SRVACQFAIL (13855L)
value ERROR_IPSEC_IKE_SRVQUERYCRED (13856L)
value ERROR_IPSEC_IKE_STRONG_CRED_AUTHORIZATION_AND_CERTMAP_FAILURE (13908L)
value ERROR_IPSEC_IKE_STRONG_CRED_AUTHORIZATION_FAILURE (13906L)
value ERROR_IPSEC_IKE_TIMED_OUT (13805L)
value ERROR_IPSEC_IKE_TOO_MANY_FILTERS (13896L)
value ERROR_IPSEC_IKE_UNEXPECTED_MESSAGE_ID (13888L)
value ERROR_IPSEC_IKE_UNKNOWN_DOI (13862L)
value ERROR_IPSEC_IKE_UNSUPPORTED_ID (13869L)
value ERROR_IPSEC_INTEGRITY_CHECK_FAILED (13915L)
value ERROR_IPSEC_INVALID_PACKET (13914L)
value ERROR_IPSEC_KEY_MODULE_IMPERSONATION_NEGOTIATION_PENDING (13901L)
value ERROR_IPSEC_MM_AUTH_EXISTS (13010L)
value ERROR_IPSEC_MM_AUTH_IN_USE (13012L)
value ERROR_IPSEC_MM_AUTH_NOT_FOUND (13011L)
value ERROR_IPSEC_MM_AUTH_PENDING_DELETION (13022L)
value ERROR_IPSEC_MM_FILTER_EXISTS (13006L)
value ERROR_IPSEC_MM_FILTER_NOT_FOUND (13007L)
value ERROR_IPSEC_MM_FILTER_PENDING_DELETION (13018L)
value ERROR_IPSEC_MM_POLICY_EXISTS (13003L)
value ERROR_IPSEC_MM_POLICY_IN_USE (13005L)
value ERROR_IPSEC_MM_POLICY_NOT_FOUND (13004L)
value ERROR_IPSEC_MM_POLICY_PENDING_DELETION (13021L)
value ERROR_IPSEC_QM_POLICY_EXISTS (13000L)
value ERROR_IPSEC_QM_POLICY_IN_USE (13002L)
value ERROR_IPSEC_QM_POLICY_NOT_FOUND (13001L)
value ERROR_IPSEC_QM_POLICY_PENDING_DELETION (13023L)
value ERROR_IPSEC_REPLAY_CHECK_FAILED (13913L)
value ERROR_IPSEC_SA_LIFETIME_EXPIRED (13911L)
value ERROR_IPSEC_THROTTLE_DROP (13918L)
value ERROR_IPSEC_TRANSPORT_FILTER_EXISTS (13008L)
value ERROR_IPSEC_TRANSPORT_FILTER_NOT_FOUND (13009L)
value ERROR_IPSEC_TRANSPORT_FILTER_PENDING_DELETION (13019L)
value ERROR_IPSEC_TUNNEL_FILTER_EXISTS (13016L)
value ERROR_IPSEC_TUNNEL_FILTER_NOT_FOUND (13017L)
value ERROR_IPSEC_TUNNEL_FILTER_PENDING_DELETION (13020L)
value ERROR_IPSEC_WRONG_SA (13912L)
value ERROR_IRQ_BUSY (1119L)
value ERROR_IS_JOINED (134L)
value ERROR_IS_JOIN_PATH (147L)
value ERROR_IS_JOIN_TARGET (133L)
value ERROR_IS_SUBSTED (135L)
value ERROR_IS_SUBST_PATH (146L)
value ERROR_IS_SUBST_TARGET (149L)
value ERROR_JOB_NO_CONTAINER (1505L)
value ERROR_JOIN_TO_JOIN (138L)
value ERROR_JOIN_TO_SUBST (140L)
value ERROR_JOURNAL_DELETE_IN_PROGRESS (1178L)
value ERROR_JOURNAL_ENTRY_DELETED (1181L)
value ERROR_JOURNAL_HOOK_SET (1430L)
value ERROR_JOURNAL_NOT_ACTIVE (1179L)
value ERROR_KERNEL_APC (738L)
value ERROR_KEY_DELETED (1018L)
value ERROR_KEY_HAS_CHILDREN (1020L)
value ERROR_KM_DRIVER_BLOCKED (1930L)
value ERROR_LABEL_TOO_LONG (154L)
value ERROR_LAST_ADMIN (1322L)
value ERROR_LB_WITHOUT_TABSTOPS (1434L)
value ERROR_LIBRARY_FULL (4322L)
value ERROR_LIBRARY_OFFLINE (4305L)
value ERROR_LICENSE_QUOTA_EXCEEDED (1395L)
value ERROR_LINUX_SUBSYSTEM_NOT_PRESENT (414L)
value ERROR_LINUX_SUBSYSTEM_UPDATE_REQUIRED (444L)
value ERROR_LISTBOX_ID_NOT_FOUND (1416L)
value ERROR_LM_CROSS_ENCRYPTION_REQUIRED (1390L)
value ERROR_LOCAL_POLICY_MODIFICATION_NOT_SUPPORTED (8653L)
value ERROR_LOCAL_USER_SESSION_KEY (1303L)
value ERROR_LOCKED (212L)
value ERROR_LOCK_FAILED (167L)
value ERROR_LOCK_VIOLATION (33L)
value ERROR_LOGIN_TIME_RESTRICTION (1239L)
value ERROR_LOGIN_WKSTA_RESTRICTION (1240L)
value ERROR_LOGON_FAILURE (1326L)
value ERROR_LOGON_NOT_GRANTED (1380L)
value ERROR_LOGON_SERVER_CONFLICT (568L)
value ERROR_LOGON_SESSION_COLLISION (1366L)
value ERROR_LOGON_SESSION_EXISTS (1363L)
value ERROR_LOGON_TYPE_NOT_GRANTED (1385L)
value ERROR_LOG_APPENDED_FLUSH_FAILED (6647L)
value ERROR_LOG_ARCHIVE_IN_PROGRESS (6633L)
value ERROR_LOG_ARCHIVE_NOT_IN_PROGRESS (6632L)
value ERROR_LOG_BLOCKS_EXHAUSTED (6605L)
value ERROR_LOG_BLOCK_INCOMPLETE (6603L)
value ERROR_LOG_BLOCK_INVALID (6609L)
value ERROR_LOG_BLOCK_VERSION (6608L)
value ERROR_LOG_CANT_DELETE (6616L)
value ERROR_LOG_CLIENT_ALREADY_REGISTERED (6636L)
value ERROR_LOG_CLIENT_NOT_REGISTERED (6637L)
value ERROR_LOG_CONTAINER_LIMIT_EXCEEDED (6617L)
value ERROR_LOG_CONTAINER_OPEN_FAILED (6641L)
value ERROR_LOG_CONTAINER_READ_FAILED (6639L)
value ERROR_LOG_CONTAINER_STATE_INVALID (6642L)
value ERROR_LOG_CONTAINER_WRITE_FAILED (6640L)
value ERROR_LOG_CORRUPTION_DETECTED (6817L)
value ERROR_LOG_DEDICATED (6631L)
value ERROR_LOG_EPHEMERAL (6634L)
value ERROR_LOG_FILE_FULL (1502L)
value ERROR_LOG_FULL (6628L)
value ERROR_LOG_FULL_HANDLER_IN_PROGRESS (6638L)
value ERROR_LOG_GROWTH_FAILED (6833L)
value ERROR_LOG_HARD_ERROR (718L)
value ERROR_LOG_INCONSISTENT_SECURITY (6646L)
value ERROR_LOG_INVALID_RANGE (6604L)
value ERROR_LOG_METADATA_CORRUPT (6612L)
value ERROR_LOG_METADATA_FLUSH_FAILED (6645L)
value ERROR_LOG_METADATA_INCONSISTENT (6614L)
value ERROR_LOG_METADATA_INVALID (6613L)
value ERROR_LOG_MULTIPLEXED (6630L)
value ERROR_LOG_NOT_ENOUGH_CONTAINERS (6635L)
value ERROR_LOG_NO_RESTART (6611L)
value ERROR_LOG_PINNED (6644L)
value ERROR_LOG_PINNED_ARCHIVE_TAIL (6623L)
value ERROR_LOG_PINNED_RESERVATION (6648L)
value ERROR_LOG_POLICY_ALREADY_INSTALLED (6619L)
value ERROR_LOG_POLICY_CONFLICT (6622L)
value ERROR_LOG_POLICY_INVALID (6621L)
value ERROR_LOG_POLICY_NOT_INSTALLED (6620L)
value ERROR_LOG_READ_CONTEXT_INVALID (6606L)
value ERROR_LOG_READ_MODE_INVALID (6610L)
value ERROR_LOG_RECORDS_RESERVED_INVALID (6625L)
value ERROR_LOG_RECORD_NONEXISTENT (6624L)
value ERROR_LOG_RESERVATION_INVALID (6615L)
value ERROR_LOG_RESIZE_INVALID_SIZE (6806L)
value ERROR_LOG_RESTART_INVALID (6607L)
value ERROR_LOG_SECTOR_INVALID (6600L)
value ERROR_LOG_SECTOR_PARITY_INVALID (6601L)
value ERROR_LOG_SECTOR_REMAPPED (6602L)
value ERROR_LOG_SPACE_RESERVED_INVALID (6626L)
value ERROR_LOG_START_OF_LOG (6618L)
value ERROR_LOG_STATE_INVALID (6643L)
value ERROR_LOG_TAIL_INVALID (6627L)
value ERROR_LONGJUMP (682L)
value ERROR_LOST_MODE_LOGON_RESTRICTION (1939L)
value ERROR_LOST_WRITEBEHIND_DATA (596L)
value ERROR_LOST_WRITEBEHIND_DATA_LOCAL_DISK_ERROR (790L)
value ERROR_LOST_WRITEBEHIND_DATA_NETWORK_DISCONNECTED (788L)
value ERROR_LOST_WRITEBEHIND_DATA_NETWORK_SERVER_ERROR (789L)
value ERROR_LUIDS_EXHAUSTED (1334L)
value ERROR_MACHINE_LOCKED (1271L)
value ERROR_MACHINE_SCOPE_NOT_ALLOWED (15666L)
value ERROR_MAGAZINE_NOT_PRESENT (1163L)
value ERROR_MALFORMED_SUBSTITUTION_STRING (14094L)
value ERROR_MAPPED_ALIGNMENT (1132L)
value ERROR_MARKED_TO_DISALLOW_WRITES (348L)
value ERROR_MARSHALL_OVERFLOW (603L)
value ERROR_MAX_SESSIONS_REACHED (353L)
value ERROR_MAX_THRDS_REACHED (164L)
value ERROR_MCA_EXCEPTION (784L)
value ERROR_MCA_INTERNAL_ERROR (15205L)
value ERROR_MCA_INVALID_CAPABILITIES_STRING (15200L)
value ERROR_MCA_INVALID_TECHNOLOGY_TYPE_RETURNED (15206L)
value ERROR_MCA_INVALID_VCP_VERSION (15201L)
value ERROR_MCA_MCCS_VERSION_MISMATCH (15203L)
value ERROR_MCA_MONITOR_VIOLATES_MCCS_SPECIFICATION (15202L)
value ERROR_MCA_OCCURED (651L)
value ERROR_MCA_UNSUPPORTED_COLOR_TEMPERATURE (15207L)
value ERROR_MCA_UNSUPPORTED_MCCS_VERSION (15204L)
value ERROR_MEDIA_CHANGED (1110L)
value ERROR_MEDIA_CHECK (679L)
value ERROR_MEDIA_INCOMPATIBLE (4315L)
value ERROR_MEDIA_NOT_AVAILABLE (4318L)
value ERROR_MEDIA_OFFLINE (4304L)
value ERROR_MEDIA_UNAVAILABLE (4308L)
value ERROR_MEDIUM_NOT_ACCESSIBLE (4323L)
value ERROR_MEMBERS_PRIMARY_GROUP (1374L)
value ERROR_MEMBER_IN_ALIAS (1378L)
value ERROR_MEMBER_IN_GROUP (1320L)
value ERROR_MEMBER_NOT_IN_ALIAS (1377L)
value ERROR_MEMBER_NOT_IN_GROUP (1321L)
value ERROR_MEMORY_HARDWARE (779L)
value ERROR_MENU_ITEM_NOT_FOUND (1456L)
value ERROR_MESSAGE_EXCEEDS_MAX_SIZE (4336L)
value ERROR_MESSAGE_SYNC_ONLY (1159L)
value ERROR_METAFILE_NOT_SUPPORTED (2003L)
value ERROR_META_EXPANSION_TOO_LONG (208L)
value ERROR_MINIVERSION_INACCESSIBLE_FROM_SPECIFIED_TRANSACTION (6810L)
value ERROR_MISSING_SYSTEMFILE (573L)
value ERROR_MOD_NOT_FOUND (126L)
value ERROR_MORE_DATA (234L)
value ERROR_MORE_WRITES (1120L)
value ERROR_MOUNT_POINT_NOT_RESOLVED (649L)
value ERROR_MP_PROCESSOR_MISMATCH (725L)
value ERROR_MRM_AUTOMERGE_ENABLED (15139L)
value ERROR_MRM_DIRECT_REF_TO_NON_DEFAULT_RESOURCE (15146L)
value ERROR_MRM_DUPLICATE_ENTRY (15119L)
value ERROR_MRM_DUPLICATE_MAP_NAME (15118L)
value ERROR_MRM_FILEPATH_TOO_LONG (15121L)
value ERROR_MRM_GENERATION_COUNT_MISMATCH (15147L)
value ERROR_MRM_INDETERMINATE_QUALIFIER_VALUE (15138L)
value ERROR_MRM_INVALID_FILE_TYPE (15112L)
value ERROR_MRM_INVALID_PRICONFIG (15111L)
value ERROR_MRM_INVALID_PRI_FILE (15126L)
value ERROR_MRM_INVALID_QUALIFIER_OPERATOR (15137L)
value ERROR_MRM_INVALID_QUALIFIER_VALUE (15114L)
value ERROR_MRM_INVALID_RESOURCE_IDENTIFIER (15120L)
value ERROR_MRM_MAP_NOT_FOUND (15135L)
value ERROR_MRM_MISSING_DEFAULT_LANGUAGE (15160L)
value ERROR_MRM_NAMED_RESOURCE_NOT_FOUND (15127L)
value ERROR_MRM_NO_CANDIDATE (15115L)
value ERROR_MRM_NO_CURRENT_VIEW_ON_THREAD (15143L)
value ERROR_MRM_NO_MATCH_OR_DEFAULT_CANDIDATE (15116L)
value ERROR_MRM_PACKAGE_NOT_FOUND (15159L)
value ERROR_MRM_RESOURCE_TYPE_MISMATCH (15117L)
value ERROR_MRM_RUNTIME_NO_DEFAULT_OR_NEUTRAL_RESOURCE (15110L)
value ERROR_MRM_SCOPE_ITEM_CONFLICT (15161L)
value ERROR_MRM_TOO_MANY_RESOURCES (15140L)
value ERROR_MRM_UNKNOWN_QUALIFIER (15113L)
value ERROR_MRM_UNSUPPORTED_DIRECTORY_TYPE (15122L)
value ERROR_MRM_UNSUPPORTED_FILE_TYPE_FOR_LOAD_UNLOAD_PRI_FILE (15142L)
value ERROR_MRM_UNSUPPORTED_FILE_TYPE_FOR_MERGE (15141L)
value ERROR_MRM_UNSUPPORTED_PROFILE_TYPE (15136L)
value ERROR_MR_MID_NOT_FOUND (317L)
value ERROR_MUI_FILE_NOT_FOUND (15100L)
value ERROR_MUI_FILE_NOT_LOADED (15105L)
value ERROR_MUI_INTLSETTINGS_INVALID_LOCALE_NAME (15108L)
value ERROR_MUI_INTLSETTINGS_UILANG_NOT_INSTALLED (15107L)
value ERROR_MUI_INVALID_FILE (15101L)
value ERROR_MUI_INVALID_LOCALE_NAME (15103L)
value ERROR_MUI_INVALID_RC_CONFIG (15102L)
value ERROR_MUI_INVALID_ULTIMATEFALLBACK_NAME (15104L)
value ERROR_MULTIPLE_FAULT_VIOLATION (640L)
value ERROR_MUTANT_LIMIT_EXCEEDED (587L)
value ERROR_MUTUAL_AUTH_FAILED (1397L)
value ERROR_NEEDS_REGISTRATION (15631L)
value ERROR_NEEDS_REMEDIATION (15612L)
value ERROR_NEGATIVE_SEEK (131L)
value ERROR_NESTING_NOT_ALLOWED (215L)
value ERROR_NETLOGON_NOT_STARTED (1792L)
value ERROR_NETNAME_DELETED (64L)
value ERROR_NETWORK_ACCESS_DENIED (65L)
value ERROR_NETWORK_ACCESS_DENIED_EDP (354L)
value ERROR_NETWORK_AUTHENTICATION_PROMPT_CANCELED (3024L)
value ERROR_NETWORK_BUSY (54L)
value ERROR_NETWORK_NOT_AVAILABLE (5035L)
value ERROR_NETWORK_UNREACHABLE (1231L)
value ERROR_NET_OPEN_FAILED (570L)
value ERROR_NET_WRITE_FAULT (88L)
value ERROR_NOACCESS (998L)
value ERROR_NODE_CANNOT_BE_CLUSTERED (5898L)
value ERROR_NODE_CANT_HOST_RESOURCE (5071L)
value ERROR_NODE_NOT_ACTIVE_CLUSTER_MEMBER (5980L)
value ERROR_NODE_NOT_AVAILABLE (5036L)
value ERROR_NOINTERFACE (632L)
value ERROR_NOLOGON_INTERDOMAIN_TRUST_ACCOUNT (1807L)
value ERROR_NOLOGON_SERVER_TRUST_ACCOUNT (1809L)
value ERROR_NOLOGON_WORKSTATION_TRUST_ACCOUNT (1808L)
value ERROR_NONCORE_GROUPS_FOUND (5937L)
value ERROR_NONE_MAPPED (1332L)
value ERROR_NONPAGED_SYSTEM_RESOURCES (1451L)
value ERROR_NON_ACCOUNT_SID (1257L)
value ERROR_NON_CSV_PATH (5950L)
value ERROR_NON_DOMAIN_SID (1258L)
value ERROR_NON_MDICHILD_WINDOW (1445L)
value ERROR_NOTHING_TO_TERMINATE (758L)
value ERROR_NOTIFICATION_GUID_ALREADY_DEFINED (309L)
value ERROR_NOTIFY_CLEANUP (745L)
value ERROR_NOTIFY_ENUM_DIR (1022L)
value ERROR_NOT_ALLOWED_ON_SYSTEM_FILE (313L)
value ERROR_NOT_ALL_ASSIGNED (1300L)
value ERROR_NOT_APPCONTAINER (4250L)
value ERROR_NOT_AUTHENTICATED (1244L)
value ERROR_NOT_A_CLOUD_FILE (376L)
value ERROR_NOT_A_CLOUD_SYNC_ROOT (405L)
value ERROR_NOT_A_DAX_VOLUME (420L)
value ERROR_NOT_A_REPARSE_POINT (4390L)
value ERROR_NOT_CAPABLE (775L)
value ERROR_NOT_CHILD_WINDOW (1442L)
value ERROR_NOT_CONNECTED (2250L)
value ERROR_NOT_CONTAINER (1207L)
value ERROR_NOT_DAX_MAPPABLE (421L)
value ERROR_NOT_DOS_DISK (26L)
value ERROR_NOT_EMPTY (4307L)
value ERROR_NOT_ENOUGH_MEMORY (8L)
value ERROR_NOT_ENOUGH_QUOTA (1816L)
value ERROR_NOT_ENOUGH_SERVER_MEMORY (1130L)
value ERROR_NOT_EXPORT_FORMAT (6008L)
value ERROR_NOT_FOUND (1168L)
value ERROR_NOT_GUI_PROCESS (1471L)
value ERROR_NOT_JOINED (136L)
value ERROR_NOT_LOCKED (158L)
value ERROR_NOT_LOGGED_ON (1245L)
value ERROR_NOT_LOGON_PROCESS (1362L)
value ERROR_NOT_OWNER (288L)
value ERROR_NOT_QUORUM_CAPABLE (5021L)
value ERROR_NOT_QUORUM_CLASS (5025L)
value ERROR_NOT_READY (21L)
value ERROR_NOT_READ_FROM_COPY (337L)
value ERROR_NOT_REDUNDANT_STORAGE (333L)
value ERROR_NOT_REGISTRY_FILE (1017L)
value ERROR_NOT_SAFEBOOT_SERVICE (1084L)
value ERROR_NOT_SAFE_MODE_DRIVER (646L)
value ERROR_NOT_SAME_DEVICE (17L)
value ERROR_NOT_SAME_OBJECT (1656L)
value ERROR_NOT_SNAPSHOT_VOLUME (6841L)
value ERROR_NOT_SUBSTED (137L)
value ERROR_NOT_SUPPORTED (50L)
value ERROR_NOT_SUPPORTED_IN_APPCONTAINER (4252L)
value ERROR_NOT_SUPPORTED_ON_DAX (360L)
value ERROR_NOT_SUPPORTED_ON_SBS (1254L)
value ERROR_NOT_SUPPORTED_ON_STANDARD_SERVER (8584L)
value ERROR_NOT_SUPPORTED_WITH_AUDITING (499L)
value ERROR_NOT_SUPPORTED_WITH_BTT (429L)
value ERROR_NOT_SUPPORTED_WITH_BYPASSIO (493L)
value ERROR_NOT_SUPPORTED_WITH_CACHED_HANDLE (509L)
value ERROR_NOT_SUPPORTED_WITH_COMPRESSION (496L)
value ERROR_NOT_SUPPORTED_WITH_DEDUPLICATION (498L)
value ERROR_NOT_SUPPORTED_WITH_ENCRYPTION (495L)
value ERROR_NOT_SUPPORTED_WITH_MONITORING (503L)
value ERROR_NOT_SUPPORTED_WITH_REPLICATION (497L)
value ERROR_NOT_SUPPORTED_WITH_SNAPSHOT (504L)
value ERROR_NOT_SUPPORTED_WITH_VIRTUALIZATION (505L)
value ERROR_NOT_TINY_STREAM (598L)
value ERROR_NO_ACE_CONDITION (804L)
value ERROR_NO_ADMIN_ACCESS_POINT (5090L)
value ERROR_NO_ASSOCIATION (1155L)
value ERROR_NO_BROWSER_SERVERS_FOUND (6118L)
value ERROR_NO_BYPASSIO_DRIVER_SUPPORT (494L)
value ERROR_NO_CALLBACK_ACTIVE (614L)
value ERROR_NO_DATA (232L)
value ERROR_NO_DATA_DETECTED (1104L)
value ERROR_NO_EFS (6004L)
value ERROR_NO_EVENT_PAIR (580L)
value ERROR_NO_GUID_TRANSLATION (560L)
value ERROR_NO_IMPERSONATION_TOKEN (1309L)
value ERROR_NO_INHERITANCE (1391L)
value ERROR_NO_LINK_TRACKING_IN_TRANSACTION (6852L)
value ERROR_NO_LOGON_SERVERS (1311L)
value ERROR_NO_LOG_SPACE (1019L)
value ERROR_NO_MATCH (1169L)
value ERROR_NO_MEDIA_IN_DRIVE (1112L)
value ERROR_NO_MORE_DEVICES (1248L)
value ERROR_NO_MORE_FILES (18L)
value ERROR_NO_MORE_ITEMS (259L)
value ERROR_NO_MORE_MATCHES (626L)
value ERROR_NO_MORE_SEARCH_HANDLES (113L)
value ERROR_NO_MORE_USER_HANDLES (1158L)
value ERROR_NO_NETWORK (1222L)
value ERROR_NO_NET_OR_BAD_PATH (1203L)
value ERROR_NO_NVRAM_RESOURCES (1470L)
value ERROR_NO_PAGEFILE (578L)
value ERROR_NO_PHYSICALLY_ALIGNED_FREE_SPACE_FOUND (408L)
value ERROR_NO_PROC_SLOTS (89L)
value ERROR_NO_PROMOTION_ACTIVE (8222L)
value ERROR_NO_QUOTAS_FOR_ACCOUNT (1302L)
value ERROR_NO_RANGES_PROCESSED (312L)
value ERROR_NO_RECOVERY_POLICY (6003L)
value ERROR_NO_RECOVERY_PROGRAM (1082L)
value ERROR_NO_SAVEPOINT_WITH_OPEN_FILES (6842L)
value ERROR_NO_SCROLLBARS (1447L)
value ERROR_NO_SECRETS (8620L)
value ERROR_NO_SECURITY_ON_OBJECT (1350L)
value ERROR_NO_SHUTDOWN_IN_PROGRESS (1116L)
value ERROR_NO_SIGNAL_SENT (205L)
value ERROR_NO_SITENAME (1919L)
value ERROR_NO_SITE_SETTINGS_OBJECT (8619L)
value ERROR_NO_SPOOL_SPACE (62L)
value ERROR_NO_SUCH_ALIAS (1376L)
value ERROR_NO_SUCH_DEVICE (433L)
value ERROR_NO_SUCH_DOMAIN (1355L)
value ERROR_NO_SUCH_GROUP (1319L)
value ERROR_NO_SUCH_LOGON_SESSION (1312L)
value ERROR_NO_SUCH_MEMBER (1387L)
value ERROR_NO_SUCH_PACKAGE (1364L)
value ERROR_NO_SUCH_PRIVILEGE (1313L)
value ERROR_NO_SUCH_SITE (1249L)
value ERROR_NO_SUCH_USER (1317L)
value ERROR_NO_SUPPORTING_DRIVES (4339L)
value ERROR_NO_SYSTEM_MENU (1437L)
value ERROR_NO_SYSTEM_RESOURCES (1450L)
value ERROR_NO_TASK_QUEUE (427L)
value ERROR_NO_TOKEN (1008L)
value ERROR_NO_TRACKING_SERVICE (1172L)
value ERROR_NO_TRUST_LSA_SECRET (1786L)
value ERROR_NO_TRUST_SAM_ACCOUNT (1787L)
value ERROR_NO_TXF_METADATA (6816L)
value ERROR_NO_UNICODE_TRANSLATION (1113L)
value ERROR_NO_USER_KEYS (6006L)
value ERROR_NO_USER_SESSION_KEY (1394L)
value ERROR_NO_VOLUME_ID (1173L)
value ERROR_NO_VOLUME_LABEL (125L)
value ERROR_NO_WILDCARD_CHARACTERS (1417L)
value ERROR_NO_WORK_DONE (235L)
value ERROR_NO_WRITABLE_DC_FOUND (8621L)
value ERROR_NO_YIELD_PERFORMED (721L)
value ERROR_NTLM_BLOCKED (1937L)
value ERROR_NT_CROSS_ENCRYPTION_REQUIRED (1386L)
value ERROR_NULL_LM_PASSWORD (1304L)
value ERROR_OBJECT_ALREADY_EXISTS (5010L)
value ERROR_OBJECT_IN_LIST (5011L)
value ERROR_OBJECT_IS_IMMUTABLE (4449L)
value ERROR_OBJECT_NAME_EXISTS (698L)
value ERROR_OBJECT_NOT_EXTERNALLY_BACKED (342L)
value ERROR_OBJECT_NOT_FOUND (4312L)
value ERROR_OBJECT_NO_LONGER_EXISTS (6807L)
value ERROR_OFFLOAD_READ_FILE_NOT_SUPPORTED (4442L)
value ERROR_OFFLOAD_READ_FLT_NOT_SUPPORTED (4440L)
value ERROR_OFFLOAD_WRITE_FILE_NOT_SUPPORTED (4443L)
value ERROR_OFFLOAD_WRITE_FLT_NOT_SUPPORTED (4441L)
value ERROR_OFFSET_ALIGNMENT_VIOLATION (327L)
value ERROR_OLD_WIN_VERSION (1150L)
value ERROR_ONLY_IF_CONNECTED (1251L)
value ERROR_OPEN_FAILED (110L)
value ERROR_OPEN_FILES (2401L)
value ERROR_OPERATION_ABORTED (995L)
value ERROR_OPERATION_IN_PROGRESS (329L)
value ERROR_OPERATION_NOT_ALLOWED_FROM_SYSTEM_COMPONENT (15145L)
value ERROR_OPERATION_NOT_SUPPORTED_IN_TRANSACTION (6853L)
value ERROR_OPLOCK_BREAK_IN_PROGRESS (742L)
value ERROR_OPLOCK_HANDLE_CLOSED (803L)
value ERROR_OPLOCK_NOT_GRANTED (300L)
value ERROR_OPLOCK_SWITCHED_TO_NEW_HANDLE (800L)
value ERROR_ORPHAN_NAME_EXHAUSTED (799L)
value ERROR_OUTOFMEMORY (14L)
value ERROR_OUT_OF_PAPER (28L)
value ERROR_OUT_OF_STRUCTURES (84L)
value ERROR_OVERRIDE_NOCHANGES (1252L)
value ERROR_PACKAGED_SERVICE_REQUIRES_ADMIN_PRIVILEGES (15656L)
value ERROR_PACKAGES_IN_USE (15618L)
value ERROR_PACKAGES_REPUTATION_CHECK_FAILED (15643L)
value ERROR_PACKAGES_REPUTATION_CHECK_TIMEDOUT (15644L)
value ERROR_PACKAGE_ALREADY_EXISTS (15611L)
value ERROR_PACKAGE_EXTERNAL_LOCATION_NOT_ALLOWED (15662L)
value ERROR_PACKAGE_LACKS_CAPABILITY_FOR_MANDATORY_STARTUPTASKS (15664L)
value ERROR_PACKAGE_LACKS_CAPABILITY_TO_DEPLOY_ON_HOST (15658L)
value ERROR_PACKAGE_MOVE_BLOCKED_BY_STREAMING (15636L)
value ERROR_PACKAGE_MOVE_FAILED (15627L)
value ERROR_PACKAGE_NAME_MISMATCH (15670L)
value ERROR_PACKAGE_NOT_REGISTERED_FOR_USER (15669L)
value ERROR_PACKAGE_NOT_SUPPORTED_ON_FILESYSTEM (15635L)
value ERROR_PACKAGE_REPOSITORY_CORRUPTED (15614L)
value ERROR_PACKAGE_STAGING_ONHOLD (15638L)
value ERROR_PACKAGE_UPDATING (15616L)
value ERROR_PAGED_SYSTEM_RESOURCES (1452L)
value ERROR_PAGEFILE_CREATE_FAILED (576L)
value ERROR_PAGEFILE_NOT_SUPPORTED (491L)
value ERROR_PAGEFILE_QUOTA (1454L)
value ERROR_PAGEFILE_QUOTA_EXCEEDED (567L)
value ERROR_PAGE_FAULT_COPY_ON_WRITE (749L)
value ERROR_PAGE_FAULT_DEMAND_ZERO (748L)
value ERROR_PAGE_FAULT_GUARD_PAGE (750L)
value ERROR_PAGE_FAULT_PAGING_FILE (751L)
value ERROR_PAGE_FAULT_TRANSITION (747L)
value ERROR_PARAMETER_QUOTA_EXCEEDED (1283L)
value ERROR_PARTIAL_COPY (299L)
value ERROR_PARTITION_FAILURE (1105L)
value ERROR_PARTITION_TERMINATING (1184L)
value ERROR_PASSWORD_CHANGE_REQUIRED (1938L)
value ERROR_PASSWORD_EXPIRED (1330L)
value ERROR_PASSWORD_MUST_CHANGE (1907L)
value ERROR_PASSWORD_RESTRICTION (1325L)
value ERROR_PATCH_MANAGED_ADVERTISED_PRODUCT (1651L)
value ERROR_PATCH_NO_SEQUENCE (1648L)
value ERROR_PATCH_PACKAGE_INVALID (1636L)
value ERROR_PATCH_PACKAGE_OPEN_FAILED (1635L)
value ERROR_PATCH_PACKAGE_REJECTED (1643L)
value ERROR_PATCH_PACKAGE_UNSUPPORTED (1637L)
value ERROR_PATCH_REMOVAL_DISALLOWED (1649L)
value ERROR_PATCH_REMOVAL_UNSUPPORTED (1646L)
value ERROR_PATCH_TARGET_NOT_FOUND (1642L)
value ERROR_PATH_BUSY (148L)
value ERROR_PATH_NOT_FOUND (3L)
value ERROR_PER_USER_TRUST_QUOTA_EXCEEDED (1932L)
value ERROR_PIPE_BUSY (231L)
value ERROR_PIPE_CONNECTED (535L)
value ERROR_PIPE_LISTENING (536L)
value ERROR_PIPE_LOCAL (229L)
value ERROR_PIPE_NOT_CONNECTED (233L)
value ERROR_PKINIT_FAILURE (1263L)
value ERROR_PLATFORM_MANIFEST_BINARY_ID_NOT_FOUND (4574L)
value ERROR_PLATFORM_MANIFEST_CATALOG_NOT_AUTHORIZED (4573L)
value ERROR_PLATFORM_MANIFEST_FILE_NOT_AUTHORIZED (4572L)
value ERROR_PLATFORM_MANIFEST_INVALID (4571L)
value ERROR_PLATFORM_MANIFEST_NOT_ACTIVE (4575L)
value ERROR_PLATFORM_MANIFEST_NOT_AUTHORIZED (4570L)
value ERROR_PLATFORM_MANIFEST_NOT_SIGNED (4576L)
value ERROR_PLUGPLAY_QUERY_VETOED (683L)
value ERROR_PNP_BAD_MPS_TABLE (671L)
value ERROR_PNP_INVALID_ID (674L)
value ERROR_PNP_IRQ_TRANSLATION_FAILED (673L)
value ERROR_PNP_QUERY_REMOVE_DEVICE_TIMEOUT (480L)
value ERROR_PNP_QUERY_REMOVE_RELATED_DEVICE_TIMEOUT (481L)
value ERROR_PNP_QUERY_REMOVE_UNRELATED_DEVICE_TIMEOUT (482L)
value ERROR_PNP_REBOOT_REQUIRED (638L)
value ERROR_PNP_RESTART_ENUMERATION (636L)
value ERROR_PNP_TRANSLATION_FAILED (672L)
value ERROR_POINT_NOT_FOUND (1171L)
value ERROR_POLICY_OBJECT_NOT_FOUND (8219L)
value ERROR_POLICY_ONLY_IN_DS (8220L)
value ERROR_POPUP_ALREADY_ACTIVE (1446L)
value ERROR_PORT_MESSAGE_TOO_LONG (546L)
value ERROR_PORT_NOT_SET (642L)
value ERROR_PORT_UNREACHABLE (1234L)
value ERROR_POSSIBLE_DEADLOCK (1131L)
value ERROR_POTENTIAL_FILE_FOUND (1180L)
value ERROR_PREDEFINED_HANDLE (714L)
value ERROR_PRIMARY_TRANSPORT_CONNECT_FAILED (746L)
value ERROR_PRINTER_ALREADY_EXISTS (1802L)
value ERROR_PRINTER_DELETED (1905L)
value ERROR_PRINTER_DRIVER_ALREADY_INSTALLED (1795L)
value ERROR_PRINTER_DRIVER_BLOCKED (3014L)
value ERROR_PRINTER_DRIVER_DOWNLOAD_NEEDED (3019L)
value ERROR_PRINTER_DRIVER_IN_USE (3001L)
value ERROR_PRINTER_DRIVER_PACKAGE_IN_USE (3015L)
value ERROR_PRINTER_DRIVER_WARNED (3013L)
value ERROR_PRINTER_HAS_JOBS_QUEUED (3009L)
value ERROR_PRINTER_NOT_FOUND (3012L)
value ERROR_PRINTER_NOT_SHAREABLE (3022L)
value ERROR_PRINTQ_FULL (61L)
value ERROR_PRINT_CANCELLED (63L)
value ERROR_PRINT_JOB_RESTART_REQUIRED (3020L)
value ERROR_PRINT_MONITOR_ALREADY_INSTALLED (3006L)
value ERROR_PRINT_MONITOR_IN_USE (3008L)
value ERROR_PRINT_PROCESSOR_ALREADY_INSTALLED (3005L)
value ERROR_PRIVATE_DIALOG_INDEX (1415L)
value ERROR_PRIVILEGE_NOT_HELD (1314L)
value ERROR_PRI_MERGE_ADD_FILE_FAILED (15151L)
value ERROR_PRI_MERGE_BUNDLE_PACKAGES_NOT_ALLOWED (15155L)
value ERROR_PRI_MERGE_INVALID_FILE_NAME (15158L)
value ERROR_PRI_MERGE_LOAD_FILE_FAILED (15150L)
value ERROR_PRI_MERGE_MAIN_PACKAGE_REQUIRED (15156L)
value ERROR_PRI_MERGE_MISSING_SCHEMA (15149L)
value ERROR_PRI_MERGE_MULTIPLE_MAIN_PACKAGES_NOT_ALLOWED (15154L)
value ERROR_PRI_MERGE_MULTIPLE_PACKAGE_FAMILIES_NOT_ALLOWED (15153L)
value ERROR_PRI_MERGE_RESOURCE_PACKAGE_REQUIRED (15157L)
value ERROR_PRI_MERGE_VERSION_MISMATCH (15148L)
value ERROR_PRI_MERGE_WRITE_FILE_FAILED (15152L)
value ERROR_PROCESS_ABORTED (1067L)
value ERROR_PROCESS_IN_JOB (760L)
value ERROR_PROCESS_IS_PROTECTED (1293L)
value ERROR_PROCESS_MODE_ALREADY_BACKGROUND (402L)
value ERROR_PROCESS_MODE_NOT_BACKGROUND (403L)
value ERROR_PROCESS_NOT_IN_JOB (759L)
value ERROR_PROC_NOT_FOUND (127L)
value ERROR_PRODUCT_UNINSTALLED (1614L)
value ERROR_PRODUCT_VERSION (1638L)
value ERROR_PROFILE_DOES_NOT_MATCH_DEVICE (2023L)
value ERROR_PROFILE_NOT_ASSOCIATED_WITH_DEVICE (2015L)
value ERROR_PROFILE_NOT_FOUND (2016L)
value ERROR_PROFILING_AT_LIMIT (553L)
value ERROR_PROFILING_NOT_STARTED (550L)
value ERROR_PROFILING_NOT_STOPPED (551L)
value ERROR_PROMOTION_ACTIVE (8221L)
value ERROR_PROTOCOL_UNREACHABLE (1233L)
value ERROR_PROVISION_OPTIONAL_PACKAGE_REQUIRES_MAIN_PACKAGE_PROVISIONED (15642L)
value ERROR_PWD_HISTORY_CONFLICT (617L)
value ERROR_PWD_TOO_LONG (657L)
value ERROR_PWD_TOO_RECENT (616L)
value ERROR_PWD_TOO_SHORT (615L)
value ERROR_QUORUMLOG_OPEN_FAILED (5028L)
value ERROR_QUORUM_DISK_NOT_FOUND (5086L)
value ERROR_QUORUM_NOT_ALLOWED_IN_THIS_GROUP (5928L)
value ERROR_QUORUM_OWNER_ALIVE (5034L)
value ERROR_QUORUM_RESOURCE (5020L)
value ERROR_QUORUM_RESOURCE_ONLINE_FAILED (5027L)
value ERROR_QUOTA_ACTIVITY (810L)
value ERROR_QUOTA_LIST_INCONSISTENT (621L)
value ERROR_RANGE_LIST_CONFLICT (627L)
value ERROR_RANGE_NOT_FOUND (644L)
value ERROR_RDP_PROTOCOL_ERROR (7065L)
value ERROR_READ_FAULT (30L)
value ERROR_RECEIVE_EXPEDITED (708L)
value ERROR_RECEIVE_PARTIAL (707L)
value ERROR_RECEIVE_PARTIAL_EXPEDITED (709L)
value ERROR_RECOVERY_FAILURE (1279L)
value ERROR_RECOVERY_FILE_CORRUPT (15619L)
value ERROR_RECOVERY_NOT_NEEDED (6821L)
value ERROR_REC_NON_EXISTENT (4005L)
value ERROR_REDIRECTION_TO_DEFAULT_ACCOUNT_NOT_ALLOWED (15657L)
value ERROR_REDIRECTOR_HAS_OPEN_HANDLES (1794L)
value ERROR_REDIR_PAUSED (72L)
value ERROR_REGISTRATION_FROM_REMOTE_DRIVE_NOT_SUPPORTED (15647L)
value ERROR_REGISTRY_CORRUPT (1015L)
value ERROR_REGISTRY_HIVE_RECOVERED (685L)
value ERROR_REGISTRY_IO_FAILED (1016L)
value ERROR_REGISTRY_QUOTA_LIMIT (613L)
value ERROR_REGISTRY_RECOVERED (1014L)
value ERROR_REG_NAT_CONSUMPTION (1261L)
value ERROR_RELOC_CHAIN_XEEDS_SEGLIM (201L)
value ERROR_REMOTE_FILE_VERSION_MISMATCH (6814L)
value ERROR_REMOTE_PRINT_CONNECTIONS_BLOCKED (1936L)
value ERROR_REMOTE_SESSION_LIMIT_EXCEEDED (1220L)
value ERROR_REMOTE_STORAGE_MEDIA_ERROR (4352L)
value ERROR_REMOTE_STORAGE_NOT_ACTIVE (4351L)
value ERROR_REMOVE_FAILED (15610L)
value ERROR_REM_NOT_LIST (51L)
value ERROR_REPARSE (741L)
value ERROR_REPARSE_ATTRIBUTE_CONFLICT (4391L)
value ERROR_REPARSE_OBJECT (755L)
value ERROR_REPARSE_POINT_ENCOUNTERED (4395L)
value ERROR_REPARSE_TAG_INVALID (4393L)
value ERROR_REPARSE_TAG_MISMATCH (4394L)
value ERROR_REPLY_MESSAGE_MISMATCH (595L)
value ERROR_REQUEST_ABORTED (1235L)
value ERROR_REQUEST_OUT_OF_SEQUENCE (776L)
value ERROR_REQUEST_PAUSED (3050L)
value ERROR_REQUEST_REFUSED (4320L)
value ERROR_REQUIRES_INTERACTIVE_WINDOWSTATION (1459L)
value ERROR_REQ_NOT_ACCEP (71L)
value ERROR_RESIDENT_FILE_NOT_SUPPORTED (334L)
value ERROR_RESILIENCY_FILE_CORRUPT (15625L)
value ERROR_RESMON_CREATE_FAILED (5017L)
value ERROR_RESMON_INVALID_STATE (5084L)
value ERROR_RESMON_ONLINE_FAILED (5018L)
value ERROR_RESMON_SYSTEM_RESOURCES_LACKING (5956L)
value ERROR_RESOURCEMANAGER_NOT_FOUND (6716L)
value ERROR_RESOURCEMANAGER_READ_ONLY (6707L)
value ERROR_RESOURCE_CALL_TIMED_OUT (5910L)
value ERROR_RESOURCE_DATA_NOT_FOUND (1812L)
value ERROR_RESOURCE_DISABLED (4309L)
value ERROR_RESOURCE_ENUM_USER_STOP (15106L)
value ERROR_RESOURCE_FAILED (5038L)
value ERROR_RESOURCE_LANG_NOT_FOUND (1815L)
value ERROR_RESOURCE_NAME_NOT_FOUND (1814L)
value ERROR_RESOURCE_NOT_AVAILABLE (5006L)
value ERROR_RESOURCE_NOT_FOUND (5007L)
value ERROR_RESOURCE_NOT_IN_AVAILABLE_STORAGE (5965L)
value ERROR_RESOURCE_NOT_ONLINE (5004L)
value ERROR_RESOURCE_NOT_PRESENT (4316L)
value ERROR_RESOURCE_ONLINE (5019L)
value ERROR_RESOURCE_PROPERTIES_STORED (5024L)
value ERROR_RESOURCE_PROPERTY_UNCHANGEABLE (5089L)
value ERROR_RESOURCE_REQUIREMENTS_CHANGED (756L)
value ERROR_RESOURCE_TYPE_NOT_FOUND (1813L)
value ERROR_RESTART_APPLICATION (1467L)
value ERROR_RESUME_HIBERNATION (727L)
value ERROR_RETRY (1237L)
value ERROR_RETURN_ADDRESS_HIJACK_ATTEMPT (1662L)
value ERROR_REVISION_MISMATCH (1306L)
value ERROR_RMODE_APP (1153L)
value ERROR_RM_ALREADY_STARTED (6822L)
value ERROR_RM_CANNOT_BE_FROZEN_FOR_SNAPSHOT (6728L)
value ERROR_RM_DISCONNECTED (6819L)
value ERROR_RM_METADATA_CORRUPT (6802L)
value ERROR_RM_NOT_ACTIVE (6801L)
value ERROR_ROLLBACK_TIMER_EXPIRED (6829L)
value ERROR_ROWSNOTRELEASED (772L)
value ERROR_RPL_NOT_ALLOWED (4006L)
value ERROR_RUNLEVEL_SWITCH_AGENT_TIMEOUT (15403L)
value ERROR_RUNLEVEL_SWITCH_IN_PROGRESS (15404L)
value ERROR_RUNLEVEL_SWITCH_TIMEOUT (15402L)
value ERROR_RWRAW_ENCRYPTED_FILE_NOT_ENCRYPTED (410L)
value ERROR_RWRAW_ENCRYPTED_INVALID_EDATAINFO_FILEOFFSET (411L)
value ERROR_RWRAW_ENCRYPTED_INVALID_EDATAINFO_FILERANGE (412L)
value ERROR_RWRAW_ENCRYPTED_INVALID_EDATAINFO_PARAMETER (413L)
value ERROR_RXACT_COMMITTED (744L)
value ERROR_RXACT_COMMIT_FAILURE (1370L)
value ERROR_RXACT_COMMIT_NECESSARY (678L)
value ERROR_RXACT_INVALID_STATE (1369L)
value ERROR_RXACT_STATE_CREATED (701L)
value ERROR_SAME_DRIVE (143L)
value ERROR_SAM_INIT_FAILURE (8541L)
value ERROR_SCOPE_NOT_FOUND (318L)
value ERROR_SCREEN_ALREADY_LOCKED (1440L)
value ERROR_SCRUB_DATA_DISABLED (332L)
value ERROR_SECONDARY_IC_PROVIDER_NOT_REGISTERED (15321L)
value ERROR_SECRET_TOO_LONG (1382L)
value ERROR_SECTION_DIRECT_MAP_ONLY (819L)
value ERROR_SECTOR_NOT_FOUND (27L)
value ERROR_SECUREBOOT_FILE_REPLACED (4426L)
value ERROR_SECUREBOOT_INVALID_POLICY (4422L)
value ERROR_SECUREBOOT_NOT_BASE_POLICY (4434L)
value ERROR_SECUREBOOT_NOT_ENABLED (4425L)
value ERROR_SECUREBOOT_NOT_SUPPLEMENTAL_POLICY (4435L)
value ERROR_SECUREBOOT_PLATFORM_ID_MISMATCH (4430L)
value ERROR_SECUREBOOT_POLICY_MISSING_ANTIROLLBACKVERSION (4429L)
value ERROR_SECUREBOOT_POLICY_NOT_AUTHORIZED (4427L)
value ERROR_SECUREBOOT_POLICY_NOT_SIGNED (4424L)
value ERROR_SECUREBOOT_POLICY_PUBLISHER_NOT_FOUND (4423L)
value ERROR_SECUREBOOT_POLICY_ROLLBACK_DETECTED (4431L)
value ERROR_SECUREBOOT_POLICY_UNKNOWN (4428L)
value ERROR_SECUREBOOT_POLICY_UPGRADE_MISMATCH (4432L)
value ERROR_SECUREBOOT_POLICY_VIOLATION (4421L)
value ERROR_SECUREBOOT_REQUIRED_POLICY_FILE_MISSING (4433L)
value ERROR_SECUREBOOT_ROLLBACK_DETECTED (4420L)
value ERROR_SECURITY_DENIES_OPERATION (447L)
value ERROR_SECURITY_STREAM_IS_INCONSISTENT (306L)
value ERROR_SEEK (25L)
value ERROR_SEEK_ON_DEVICE (132L)
value ERROR_SEGMENT_NOTIFICATION (702L)
value ERROR_SEM_IS_SET (102L)
value ERROR_SEM_NOT_FOUND (187L)
value ERROR_SEM_OWNER_DIED (105L)
value ERROR_SEM_TIMEOUT (121L)
value ERROR_SEM_USER_LIMIT (106L)
value ERROR_SERIAL_NO_DEVICE (1118L)
value ERROR_SERVER_DISABLED (1341L)
value ERROR_SERVER_HAS_OPEN_HANDLES (1811L)
value ERROR_SERVER_NOT_DISABLED (1342L)
value ERROR_SERVER_SHUTDOWN_IN_PROGRESS (1255L)
value ERROR_SERVER_SID_MISMATCH (628L)
value ERROR_SERVER_TRANSPORT_CONFLICT (816L)
value ERROR_SERVICES_FAILED_AUTOSTART (15405L)
value ERROR_SERVICE_ALREADY_RUNNING (1056L)
value ERROR_SERVICE_CANNOT_ACCEPT_CTRL (1061L)
value ERROR_SERVICE_DATABASE_LOCKED (1055L)
value ERROR_SERVICE_DEPENDENCY_DELETED (1075L)
value ERROR_SERVICE_DEPENDENCY_FAIL (1068L)
value ERROR_SERVICE_DISABLED (1058L)
value ERROR_SERVICE_DOES_NOT_EXIST (1060L)
value ERROR_SERVICE_EXISTS (1073L)
value ERROR_SERVICE_EXISTS_AS_NON_PACKAGED_SERVICE (15655L)
value ERROR_SERVICE_LOGON_FAILED (1069L)
value ERROR_SERVICE_MARKED_FOR_DELETE (1072L)
value ERROR_SERVICE_NEVER_STARTED (1077L)
value ERROR_SERVICE_NOTIFICATION (716L)
value ERROR_SERVICE_NOTIFY_CLIENT_LAGGING (1294L)
value ERROR_SERVICE_NOT_ACTIVE (1062L)
value ERROR_SERVICE_NOT_FOUND (1243L)
value ERROR_SERVICE_NOT_IN_EXE (1083L)
value ERROR_SERVICE_NO_THREAD (1054L)
value ERROR_SERVICE_REQUEST_TIMEOUT (1053L)
value ERROR_SERVICE_SPECIFIC_ERROR (1066L)
value ERROR_SERVICE_START_HANG (1070L)
value ERROR_SESSION_CREDENTIAL_CONFLICT (1219L)
value ERROR_SESSION_KEY_TOO_SHORT (501L)
value ERROR_SETCOUNT_ON_BAD_LB (1433L)
value ERROR_SETMARK_DETECTED (1103L)
value ERROR_SET_CONTEXT_DENIED (1660L)
value ERROR_SET_NOT_FOUND (1170L)
value ERROR_SET_POWER_STATE_FAILED (1141L)
value ERROR_SET_POWER_STATE_VETOED (1140L)
value ERROR_SHARED_POLICY (8218L)
value ERROR_SHARING_BUFFER_EXCEEDED (36L)
value ERROR_SHARING_PAUSED (70L)
value ERROR_SHARING_VIOLATION (32L)
value ERROR_SHORT_NAMES_NOT_ENABLED_ON_VOLUME (305L)
value ERROR_SHUTDOWN_CLUSTER (5008L)
value ERROR_SHUTDOWN_DISKS_NOT_IN_MAINTENANCE_MODE (1192L)
value ERROR_SHUTDOWN_IN_PROGRESS (1115L)
value ERROR_SHUTDOWN_IS_SCHEDULED (1190L)
value ERROR_SHUTDOWN_USERS_LOGGED_ON (1191L)
value ERROR_SIGNAL_PENDING (162L)
value ERROR_SIGNAL_REFUSED (156L)
value ERROR_SIGNED_PACKAGE_INVALID_PUBLISHER_NAMESPACE (15661L)
value ERROR_SINGLETON_RESOURCE_INSTALLED_IN_ACTIVE_USER (15653L)
value ERROR_SINGLE_INSTANCE_APP (1152L)
value ERROR_SMARTCARD_SUBSYSTEM_FAILURE (1264L)
value ERROR_SMB_GUEST_LOGON_BLOCKED (1272L)
value ERROR_SMI_PRIMITIVE_INSTALLER_FAILED (14108L)
value ERROR_SMR_GARBAGE_COLLECTION_REQUIRED (4445L)
value ERROR_SOME_NOT_MAPPED (1301L)
value ERROR_SOURCE_ELEMENT_EMPTY (1160L)
value ERROR_SPARSE_FILE_NOT_SUPPORTED (490L)
value ERROR_SPARSE_NOT_ALLOWED_IN_TRANSACTION (6844L)
value ERROR_SPECIAL_ACCOUNT (1371L)
value ERROR_SPECIAL_GROUP (1372L)
value ERROR_SPECIAL_USER (1373L)
value ERROR_SPL_NO_ADDJOB (3004L)
value ERROR_SPL_NO_STARTDOC (3003L)
value ERROR_SPOOL_FILE_NOT_FOUND (3002L)
value ERROR_SRC_SRV_DLL_LOAD_FAILED (428L)
value ERROR_STACK_BUFFER_OVERRUN (1282L)
value ERROR_STACK_OVERFLOW (1001L)
value ERROR_STACK_OVERFLOW_READ (599L)
value ERROR_STAGEFROMUPDATEAGENT_PACKAGE_NOT_APPLICABLE (15668L)
value ERROR_STATE_COMPOSITE_SETTING_VALUE_SIZE_LIMIT_EXCEEDED (15815L)
value ERROR_STATE_CONTAINER_NAME_SIZE_LIMIT_EXCEEDED (15818L)
value ERROR_STATE_CREATE_CONTAINER_FAILED (15805L)
value ERROR_STATE_DELETE_CONTAINER_FAILED (15806L)
value ERROR_STATE_DELETE_SETTING_FAILED (15809L)
value ERROR_STATE_ENUMERATE_CONTAINER_FAILED (15813L)
value ERROR_STATE_ENUMERATE_SETTINGS_FAILED (15814L)
value ERROR_STATE_GET_VERSION_FAILED (15801L)
value ERROR_STATE_LOAD_STORE_FAILED (15800L)
value ERROR_STATE_OPEN_CONTAINER_FAILED (15804L)
value ERROR_STATE_QUERY_SETTING_FAILED (15810L)
value ERROR_STATE_READ_COMPOSITE_SETTING_FAILED (15811L)
value ERROR_STATE_READ_SETTING_FAILED (15807L)
value ERROR_STATE_SETTING_NAME_SIZE_LIMIT_EXCEEDED (15817L)
value ERROR_STATE_SETTING_VALUE_SIZE_LIMIT_EXCEEDED (15816L)
value ERROR_STATE_SET_VERSION_FAILED (15802L)
value ERROR_STATE_STRUCTURED_RESET_FAILED (15803L)
value ERROR_STATE_WRITE_COMPOSITE_SETTING_FAILED (15812L)
value ERROR_STATE_WRITE_SETTING_FAILED (15808L)
value ERROR_STATIC_INIT (4002L)
value ERROR_STOPPED_ON_SYMLINK (681L)
value ERROR_STORAGE_LOST_DATA_PERSISTENCE (368L)
value ERROR_STORAGE_RESERVE_ALREADY_EXISTS (418L)
value ERROR_STORAGE_RESERVE_DOES_NOT_EXIST (417L)
value ERROR_STORAGE_RESERVE_ID_INVALID (416L)
value ERROR_STORAGE_RESERVE_NOT_EMPTY (419L)
value ERROR_STORAGE_STACK_ACCESS_DENIED (472L)
value ERROR_STORAGE_TOPOLOGY_ID_MISMATCH (345L)
value ERROR_STREAM_MINIVERSION_NOT_FOUND (6808L)
value ERROR_STREAM_MINIVERSION_NOT_VALID (6809L)
value ERROR_STRICT_CFG_VIOLATION (1657L)
value ERROR_SUBST_TO_JOIN (141L)
value ERROR_SUBST_TO_SUBST (139L)
value ERROR_SUCCESS (0cL)
value ERROR_SUCCESS_REBOOT_INITIATED (1641L)
value ERROR_SUCCESS_REBOOT_REQUIRED (3010L)
value ERROR_SUCCESS_RESTART_REQUIRED (3011L)
value ERROR_SWAPERROR (999L)
value ERROR_SXS_ACTIVATION_CONTEXT_DISABLED (14006L)
value ERROR_SXS_ASSEMBLY_IS_NOT_A_DEPLOYMENT (14103L)
value ERROR_SXS_ASSEMBLY_MISSING (14081L)
value ERROR_SXS_ASSEMBLY_NOT_FOUND (14003L)
value ERROR_SXS_ASSEMBLY_NOT_LOCKED (14097L)
value ERROR_SXS_CANT_GEN_ACTCTX (14001L)
value ERROR_SXS_COMPONENT_STORE_CORRUPT (14098L)
value ERROR_SXS_CORRUPTION (14083L)
value ERROR_SXS_CORRUPT_ACTIVATION_STACK (14082L)
value ERROR_SXS_DUPLICATE_ACTIVATABLE_CLASS (14111L)
value ERROR_SXS_DUPLICATE_ASSEMBLY_NAME (14027L)
value ERROR_SXS_DUPLICATE_CLSID (14023L)
value ERROR_SXS_DUPLICATE_DLL_NAME (14021L)
value ERROR_SXS_DUPLICATE_IID (14024L)
value ERROR_SXS_DUPLICATE_PROGID (14026L)
value ERROR_SXS_DUPLICATE_TLBID (14025L)
value ERROR_SXS_DUPLICATE_WINDOWCLASS_NAME (14022L)
value ERROR_SXS_EARLY_DEACTIVATION (14084L)
value ERROR_SXS_FILE_HASH_MISMATCH (14028L)
value ERROR_SXS_FILE_HASH_MISSING (14110L)
value ERROR_SXS_FILE_NOT_PART_OF_ASSEMBLY (14104L)
value ERROR_SXS_IDENTITIES_DIFFERENT (14102L)
value ERROR_SXS_IDENTITY_DUPLICATE_ATTRIBUTE (14092L)
value ERROR_SXS_IDENTITY_PARSE_ERROR (14093L)
value ERROR_SXS_INCORRECT_PUBLIC_KEY_TOKEN (14095L)
value ERROR_SXS_INVALID_ACTCTXDATA_FORMAT (14002L)
value ERROR_SXS_INVALID_ASSEMBLY_IDENTITY_ATTRIBUTE (14017L)
value ERROR_SXS_INVALID_ASSEMBLY_IDENTITY_ATTRIBUTE_NAME (14080L)
value ERROR_SXS_INVALID_DEACTIVATION (14085L)
value ERROR_SXS_INVALID_IDENTITY_ATTRIBUTE_NAME (14091L)
value ERROR_SXS_INVALID_IDENTITY_ATTRIBUTE_VALUE (14090L)
value ERROR_SXS_INVALID_XML_NAMESPACE_URI (14014L)
value ERROR_SXS_KEY_NOT_FOUND (14007L)
value ERROR_SXS_LEAF_MANIFEST_DEPENDENCY_NOT_INSTALLED (14016L)
value ERROR_SXS_MANIFEST_FORMAT_ERROR (14004L)
value ERROR_SXS_MANIFEST_IDENTITY_SAME_BUT_CONTENTS_DIFFERENT (14101L)
value ERROR_SXS_MANIFEST_INVALID_REQUIRED_DEFAULT_NAMESPACE (14019L)
value ERROR_SXS_MANIFEST_MISSING_REQUIRED_DEFAULT_NAMESPACE (14018L)
value ERROR_SXS_MANIFEST_PARSE_ERROR (14005L)
value ERROR_SXS_MANIFEST_TOO_BIG (14105L)
value ERROR_SXS_MISSING_ASSEMBLY_IDENTITY_ATTRIBUTE (14079L)
value ERROR_SXS_MULTIPLE_DEACTIVATION (14086L)
value ERROR_SXS_POLICY_PARSE_ERROR (14029L)
value ERROR_SXS_PRIVATE_MANIFEST_CROSS_PATH_WITH_REPARSE_POINT (14020L)
value ERROR_SXS_PROCESS_DEFAULT_ALREADY_SET (14011L)
value ERROR_SXS_PROCESS_TERMINATION_REQUESTED (14087L)
value ERROR_SXS_PROTECTION_CATALOG_FILE_MISSING (14078L)
value ERROR_SXS_PROTECTION_CATALOG_NOT_VALID (14076L)
value ERROR_SXS_PROTECTION_PUBLIC_KEY_TOO_SHORT (14075L)
value ERROR_SXS_PROTECTION_RECOVERY_FAILED (14074L)
value ERROR_SXS_RELEASE_ACTIVATION_CONTEXT (14088L)
value ERROR_SXS_ROOT_MANIFEST_DEPENDENCY_NOT_INSTALLED (14015L)
value ERROR_SXS_SECTION_NOT_FOUND (14000L)
value ERROR_SXS_SETTING_NOT_REGISTERED (14106L)
value ERROR_SXS_SYSTEM_DEFAULT_ACTIVATION_CONTEXT_EMPTY (14089L)
value ERROR_SXS_THREAD_QUERIES_DISABLED (14010L)
value ERROR_SXS_TRANSACTION_CLOSURE_INCOMPLETE (14107L)
value ERROR_SXS_UNKNOWN_ENCODING (14013L)
value ERROR_SXS_UNKNOWN_ENCODING_GROUP (14012L)
value ERROR_SXS_UNTRANSLATABLE_HRESULT (14077L)
value ERROR_SXS_VERSION_CONFLICT (14008L)
value ERROR_SXS_WRONG_SECTION_TYPE (14009L)
value ERROR_SXS_XML_E_BADCHARDATA (14036L)
value ERROR_SXS_XML_E_BADCHARINSTRING (14034L)
value ERROR_SXS_XML_E_BADNAMECHAR (14033L)
value ERROR_SXS_XML_E_BADPEREFINSUBSET (14059L)
value ERROR_SXS_XML_E_BADSTARTNAMECHAR (14032L)
value ERROR_SXS_XML_E_BADXMLCASE (14069L)
value ERROR_SXS_XML_E_BADXMLDECL (14056L)
value ERROR_SXS_XML_E_COMMENTSYNTAX (14031L)
value ERROR_SXS_XML_E_DUPLICATEATTRIBUTE (14053L)
value ERROR_SXS_XML_E_EXPECTINGCLOSEQUOTE (14045L)
value ERROR_SXS_XML_E_EXPECTINGTAGEND (14038L)
value ERROR_SXS_XML_E_INCOMPLETE_ENCODING (14043L)
value ERROR_SXS_XML_E_INTERNALERROR (14041L)
value ERROR_SXS_XML_E_INVALIDATROOTLEVEL (14055L)
value ERROR_SXS_XML_E_INVALIDENCODING (14067L)
value ERROR_SXS_XML_E_INVALIDSWITCH (14068L)
value ERROR_SXS_XML_E_INVALID_DECIMAL (14047L)
value ERROR_SXS_XML_E_INVALID_HEXIDECIMAL (14048L)
value ERROR_SXS_XML_E_INVALID_STANDALONE (14070L)
value ERROR_SXS_XML_E_INVALID_UNICODE (14049L)
value ERROR_SXS_XML_E_INVALID_VERSION (14072L)
value ERROR_SXS_XML_E_MISSINGEQUALS (14073L)
value ERROR_SXS_XML_E_MISSINGQUOTE (14030L)
value ERROR_SXS_XML_E_MISSINGROOT (14057L)
value ERROR_SXS_XML_E_MISSINGSEMICOLON (14039L)
value ERROR_SXS_XML_E_MISSINGWHITESPACE (14037L)
value ERROR_SXS_XML_E_MISSING_PAREN (14044L)
value ERROR_SXS_XML_E_MULTIPLEROOTS (14054L)
value ERROR_SXS_XML_E_MULTIPLE_COLONS (14046L)
value ERROR_SXS_XML_E_RESERVEDNAMESPACE (14066L)
value ERROR_SXS_XML_E_UNBALANCEDPAREN (14040L)
value ERROR_SXS_XML_E_UNCLOSEDCDATA (14065L)
value ERROR_SXS_XML_E_UNCLOSEDCOMMENT (14063L)
value ERROR_SXS_XML_E_UNCLOSEDDECL (14064L)
value ERROR_SXS_XML_E_UNCLOSEDENDTAG (14061L)
value ERROR_SXS_XML_E_UNCLOSEDSTARTTAG (14060L)
value ERROR_SXS_XML_E_UNCLOSEDSTRING (14062L)
value ERROR_SXS_XML_E_UNCLOSEDTAG (14052L)
value ERROR_SXS_XML_E_UNEXPECTEDENDTAG (14051L)
value ERROR_SXS_XML_E_UNEXPECTEDEOF (14058L)
value ERROR_SXS_XML_E_UNEXPECTED_STANDALONE (14071L)
value ERROR_SXS_XML_E_UNEXPECTED_WHITESPACE (14042L)
value ERROR_SXS_XML_E_WHITESPACEORQUESTIONMARK (14050L)
value ERROR_SXS_XML_E_XMLDECLSYNTAX (14035L)
value ERROR_SYMLINK_CLASS_DISABLED (1463L)
value ERROR_SYMLINK_NOT_SUPPORTED (1464L)
value ERROR_SYNCHRONIZATION_REQUIRED (569L)
value ERROR_SYNC_FOREGROUND_REFRESH_REQUIRED (1274L)
value ERROR_SYSTEM_DEVICE_NOT_FOUND (15299L)
value ERROR_SYSTEM_HIVE_TOO_LARGE (653L)
value ERROR_SYSTEM_IMAGE_BAD_SIGNATURE (637L)
value ERROR_SYSTEM_INTEGRITY_INVALID_POLICY (4552L)
value ERROR_SYSTEM_INTEGRITY_POLICY_NOT_SIGNED (4553L)
value ERROR_SYSTEM_INTEGRITY_POLICY_VIOLATION (4551L)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_DANGEROUS_EXT (4558L)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_MALICIOUS (4556L)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_OFFLINE (4559L)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_PUA (4557L)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_UNATTAINABLE (4581L)
value ERROR_SYSTEM_INTEGRITY_REPUTATION_UNFRIENDLY_FILE (4580L)
value ERROR_SYSTEM_INTEGRITY_ROLLBACK_DETECTED (4550L)
value ERROR_SYSTEM_INTEGRITY_SUPPLEMENTAL_POLICY_NOT_AUTHORIZED (4555L)
value ERROR_SYSTEM_INTEGRITY_TOO_MANY_POLICIES (4554L)
value ERROR_SYSTEM_NEEDS_REMEDIATION (15623L)
value ERROR_SYSTEM_POWERSTATE_COMPLEX_TRANSITION (783L)
value ERROR_SYSTEM_POWERSTATE_TRANSITION (782L)
value ERROR_SYSTEM_PROCESS_TERMINATED (591L)
value ERROR_SYSTEM_SHUTDOWN (641L)
value ERROR_SYSTEM_TRACE (150L)
value ERROR_TAG_NOT_FOUND (2012L)
value ERROR_TAG_NOT_PRESENT (2013L)
value ERROR_THREAD_ALREADY_IN_TASK (1552L)
value ERROR_THREAD_MODE_ALREADY_BACKGROUND (400L)
value ERROR_THREAD_MODE_NOT_BACKGROUND (401L)
value ERROR_THREAD_NOT_IN_PROCESS (566L)
value ERROR_THREAD_WAS_SUSPENDED (699L)
value ERROR_TIMEOUT (1460L)
value ERROR_TIMER_NOT_CANCELED (541L)
value ERROR_TIMER_RESOLUTION_NOT_SET (607L)
value ERROR_TIMER_RESUME_IGNORED (722L)
value ERROR_TIME_SENSITIVE_THREAD (422L)
value ERROR_TIME_SKEW (1398L)
value ERROR_TLW_WITH_WSCHILD (1406L)
value ERROR_TM_IDENTITY_MISMATCH (6845L)
value ERROR_TM_INITIALIZATION_FAILED (6706L)
value ERROR_TM_VOLATILE (6828L)
value ERROR_TOKEN_ALREADY_IN_USE (1375L)
value ERROR_TOO_MANY_CMDS (56L)
value ERROR_TOO_MANY_CONTEXT_IDS (1384L)
value ERROR_TOO_MANY_DESCRIPTORS (331L)
value ERROR_TOO_MANY_LINKS (1142L)
value ERROR_TOO_MANY_LUIDS_REQUESTED (1333L)
value ERROR_TOO_MANY_MODULES (214L)
value ERROR_TOO_MANY_MUXWAITERS (152L)
value ERROR_TOO_MANY_NAMES (68L)
value ERROR_TOO_MANY_OPEN_FILES (4L)
value ERROR_TOO_MANY_POSTS (298L)
value ERROR_TOO_MANY_SECRETS (1381L)
value ERROR_TOO_MANY_SEMAPHORES (100L)
value ERROR_TOO_MANY_SEM_REQUESTS (103L)
value ERROR_TOO_MANY_SESS (69L)
value ERROR_TOO_MANY_SIDS (1389L)
value ERROR_TOO_MANY_TCBS (155L)
value ERROR_TOO_MANY_THREADS (565L)
value ERROR_TRANSACTED_MAPPING_UNSUPPORTED_REMOTE (6834L)
value ERROR_TRANSACTIONAL_CONFLICT (6800L)
value ERROR_TRANSACTIONAL_OPEN_NOT_ALLOWED (6832L)
value ERROR_TRANSACTIONMANAGER_IDENTITY_MISMATCH (6727L)
value ERROR_TRANSACTIONMANAGER_NOT_FOUND (6718L)
value ERROR_TRANSACTIONMANAGER_NOT_ONLINE (6719L)
value ERROR_TRANSACTIONMANAGER_RECOVERY_NAME_COLLISION (6720L)
value ERROR_TRANSACTIONS_NOT_FROZEN (6839L)
value ERROR_TRANSACTIONS_UNSUPPORTED_REMOTE (6805L)
value ERROR_TRANSACTION_ALREADY_ABORTED (6704L)
value ERROR_TRANSACTION_ALREADY_COMMITTED (6705L)
value ERROR_TRANSACTION_FREEZE_IN_PROGRESS (6840L)
value ERROR_TRANSACTION_INTEGRITY_VIOLATED (6726L)
value ERROR_TRANSACTION_INVALID_MARSHALL_BUFFER (6713L)
value ERROR_TRANSACTION_MUST_WRITETHROUGH (6729L)
value ERROR_TRANSACTION_NOT_ACTIVE (6701L)
value ERROR_TRANSACTION_NOT_ENLISTED (6855L)
value ERROR_TRANSACTION_NOT_FOUND (6715L)
value ERROR_TRANSACTION_NOT_JOINED (6708L)
value ERROR_TRANSACTION_NOT_REQUESTED (6703L)
value ERROR_TRANSACTION_NOT_ROOT (6721L)
value ERROR_TRANSACTION_NO_SUPERIOR (6730L)
value ERROR_TRANSACTION_OBJECT_EXPIRED (6722L)
value ERROR_TRANSACTION_PROPAGATION_FAILED (6711L)
value ERROR_TRANSACTION_RECORD_TOO_LONG (6724L)
value ERROR_TRANSACTION_REQUEST_NOT_VALID (6702L)
value ERROR_TRANSACTION_REQUIRED_PROMOTION (6837L)
value ERROR_TRANSACTION_RESPONSE_NOT_ENLISTED (6723L)
value ERROR_TRANSACTION_SCOPE_CALLBACKS_NOT_SET (6836L)
value ERROR_TRANSACTION_SUPERIOR_EXISTS (6709L)
value ERROR_TRANSFORM_NOT_SUPPORTED (2004L)
value ERROR_TRANSLATION_COMPLETE (757L)
value ERROR_TRANSPORT_FULL (4328L)
value ERROR_TRUSTED_DOMAIN_FAILURE (1788L)
value ERROR_TRUSTED_RELATIONSHIP_FAILURE (1789L)
value ERROR_TRUST_FAILURE (1790L)
value ERROR_TS_INCOMPATIBLE_SESSIONS (7069L)
value ERROR_TS_VIDEO_SUBSYSTEM_ERROR (7070L)
value ERROR_TXF_ATTRIBUTE_CORRUPT (6830L)
value ERROR_TXF_DIR_NOT_EMPTY (6826L)
value ERROR_TXF_METADATA_ALREADY_PRESENT (6835L)
value ERROR_UNABLE_TO_CLEAN (4311L)
value ERROR_UNABLE_TO_EJECT_MOUNTED_MEDIA (4330L)
value ERROR_UNABLE_TO_INVENTORY_DRIVE (4325L)
value ERROR_UNABLE_TO_INVENTORY_SLOT (4326L)
value ERROR_UNABLE_TO_INVENTORY_TRANSPORT (4327L)
value ERROR_UNABLE_TO_LOAD_MEDIUM (4324L)
value ERROR_UNABLE_TO_LOCK_MEDIA (1108L)
value ERROR_UNABLE_TO_MOVE_REPLACEMENT (1176L)
value ERROR_UNABLE_TO_REMOVE_REPLACED (1175L)
value ERROR_UNABLE_TO_UNLOAD_MEDIA (1109L)
value ERROR_UNDEFINED_CHARACTER (583L)
value ERROR_UNDEFINED_SCOPE (319L)
value ERROR_UNEXPECTED_MM_CREATE_ERR (556L)
value ERROR_UNEXPECTED_MM_EXTEND_ERR (558L)
value ERROR_UNEXPECTED_MM_MAP_ERROR (557L)
value ERROR_UNEXPECTED_NTCACHEMANAGER_ERROR (443L)
value ERROR_UNEXPECTED_OMID (4334L)
value ERROR_UNEXP_NET_ERR (59L)
value ERROR_UNHANDLED_EXCEPTION (574L)
value ERROR_UNIDENTIFIED_ERROR (1287L)
value ERROR_UNKNOWN_COMPONENT (1607L)
value ERROR_UNKNOWN_FEATURE (1606L)
value ERROR_UNKNOWN_PATCH (1647L)
value ERROR_UNKNOWN_PORT (1796L)
value ERROR_UNKNOWN_PRINTER_DRIVER (1797L)
value ERROR_UNKNOWN_PRINTPROCESSOR (1798L)
value ERROR_UNKNOWN_PRINT_MONITOR (3000L)
value ERROR_UNKNOWN_PRODUCT (1605L)
value ERROR_UNKNOWN_PROPERTY (1608L)
value ERROR_UNKNOWN_REVISION (1305L)
value ERROR_UNMAPPED_SUBSTITUTION_STRING (14096L)
value ERROR_UNRECOGNIZED_MEDIA (1785L)
value ERROR_UNRECOGNIZED_VOLUME (1005L)
value ERROR_UNSATISFIED_DEPENDENCIES (441L)
value ERROR_UNSIGNED_PACKAGE_INVALID_CONTENT (15659L)
value ERROR_UNSIGNED_PACKAGE_INVALID_PUBLISHER_NAMESPACE (15660L)
value ERROR_UNSUPPORTED_COMPRESSION (618L)
value ERROR_UNSUPPORTED_TYPE (1630L)
value ERROR_UNTRUSTED_MOUNT_POINT (448L)
value ERROR_UNWIND (542L)
value ERROR_UNWIND_CONSOLIDATE (684L)
value ERROR_USER_APC (737L)
value ERROR_USER_DELETE_TRUST_QUOTA_EXCEEDED (1934L)
value ERROR_USER_EXISTS (1316L)
value ERROR_USER_MAPPED_FILE (1224L)
value ERROR_USER_PROFILE_LOAD (500L)
value ERROR_VALIDATE_CONTINUE (625L)
value ERROR_VC_DISCONNECTED (240L)
value ERROR_VDM_DISALLOWED (1286L)
value ERROR_VDM_HARD_ERROR (593L)
value ERROR_VERIFIER_STOP (537L)
value ERROR_VERSION_PARSE_ERROR (777L)
value ERROR_VIRUS_DELETED (226L)
value ERROR_VIRUS_INFECTED (225L)
value ERROR_VOLSNAP_HIBERNATE_READY (761L)
value ERROR_VOLSNAP_PREPARE_HIBERNATE (655L)
value ERROR_VOLUME_CONTAINS_SYS_FILES (4337L)
value ERROR_VOLUME_DIRTY (6851L)
value ERROR_VOLUME_MOUNTED (743L)
value ERROR_VOLUME_NOT_CLUSTER_ALIGNED (407L)
value ERROR_VOLUME_NOT_SIS_ENABLED (4500L)
value ERROR_VOLUME_NOT_SUPPORTED (492L)
value ERROR_VOLUME_NOT_SUPPORT_EFS (6014L)
value ERROR_VOLUME_WRITE_ACCESS_DENIED (508L)
value ERROR_VRF_VOLATILE_CFG_AND_IO_ENABLED (3080L)
value ERROR_VRF_VOLATILE_NMI_REGISTERED (3086L)
value ERROR_VRF_VOLATILE_NOT_RUNNABLE_SYSTEM (3083L)
value ERROR_VRF_VOLATILE_NOT_STOPPABLE (3081L)
value ERROR_VRF_VOLATILE_NOT_SUPPORTED_RULECLASS (3084L)
value ERROR_VRF_VOLATILE_PROTECTED_DRIVER (3085L)
value ERROR_VRF_VOLATILE_SAFE_MODE (3082L)
value ERROR_VRF_VOLATILE_SETTINGS_CONFLICT (3087L)
value ERROR_VSM_DMA_PROTECTION_NOT_IN_USE (4561L)
value ERROR_VSM_NOT_INITIALIZED (4560L)
value ERROR_WAIT_FOR_OPLOCK (765L)
value ERROR_WAIT_NO_CHILDREN (128L)
value ERROR_WAKE_SYSTEM (730L)
value ERROR_WAKE_SYSTEM_DEBUGGER (675L)
value ERROR_WAS_LOCKED (717L)
value ERROR_WAS_UNLOCKED (715L)
value ERROR_WEAK_WHFBKEY_BLOCKED (8651L)
value ERROR_WINDOW_NOT_COMBOBOX (1423L)
value ERROR_WINDOW_NOT_DIALOG (1420L)
value ERROR_WINDOW_OF_OTHER_THREAD (1408L)
value ERROR_WINS_INTERNAL (4000L)
value ERROR_WIP_ENCRYPTION_FAILED (6023L)
value ERROR_WMI_ALREADY_DISABLED (4212L)
value ERROR_WMI_ALREADY_ENABLED (4206L)
value ERROR_WMI_DP_FAILED (4209L)
value ERROR_WMI_DP_NOT_FOUND (4204L)
value ERROR_WMI_GUID_DISCONNECTED (4207L)
value ERROR_WMI_GUID_NOT_FOUND (4200L)
value ERROR_WMI_INSTANCE_NOT_FOUND (4201L)
value ERROR_WMI_INVALID_MOF (4210L)
value ERROR_WMI_INVALID_REGINFO (4211L)
value ERROR_WMI_ITEMID_NOT_FOUND (4202L)
value ERROR_WMI_READ_ONLY (4213L)
value ERROR_WMI_SERVER_UNAVAILABLE (4208L)
value ERROR_WMI_SET_FAILURE (4214L)
value ERROR_WMI_TRY_AGAIN (4203L)
value ERROR_WMI_UNRESOLVED_INSTANCE_REF (4205L)
value ERROR_WOF_FILE_RESOURCE_TABLE_CORRUPT (4448L)
value ERROR_WOF_WIM_HEADER_CORRUPT (4446L)
value ERROR_WOF_WIM_RESOURCE_TABLE_CORRUPT (4447L)
value ERROR_WORKING_SET_QUOTA (1453L)
value ERROR_WOW_ASSERTION (670L)
value ERROR_WRITE_FAULT (29L)
value ERROR_WRITE_PROTECT (19L)
value ERROR_WRONG_COMPARTMENT (1468L)
value ERROR_WRONG_DISK (34L)
value ERROR_WRONG_EFS (6005L)
value ERROR_WRONG_PASSWORD (1323L)
value ERROR_WRONG_TARGET_NAME (1396L)
value ERROR_XMLDSIG_ERROR (1466L)
value ERROR_XML_ENCODING_MISMATCH (14100L)
value ERROR_XML_PARSE_ERROR (1465L)
value ESB_DISABLE_LTUP (ESB_DISABLE_LEFT)
value ESB_DISABLE_RTDN (ESB_DISABLE_RIGHT)
value ESPIPE (29)
value ESRCH (3)
value ETIME (137)
value ETIMEDOUT (138)
value ETXTBSY (139)
value EVENPARITY (2)
value EVENTLOG_FULL_INFO (0)
value EWOULDBLOCK (140)
value EXCEPTION_ACCESS_VIOLATION (STATUS_ACCESS_VIOLATION)
value EXCEPTION_ARRAY_BOUNDS_EXCEEDED (STATUS_ARRAY_BOUNDS_EXCEEDED)
value EXCEPTION_BREAKPOINT (STATUS_BREAKPOINT)
value EXCEPTION_CONTINUE_SEARCH (0)
value EXCEPTION_DATATYPE_MISALIGNMENT (STATUS_DATATYPE_MISALIGNMENT)
value EXCEPTION_DEBUG_EVENT (1)
value EXCEPTION_EXECUTE_FAULT (8)
value EXCEPTION_EXECUTE_HANDLER (1)
value EXCEPTION_FLT_DENORMAL_OPERAND (STATUS_FLOAT_DENORMAL_OPERAND)
value EXCEPTION_FLT_DIVIDE_BY_ZERO (STATUS_FLOAT_DIVIDE_BY_ZERO)
value EXCEPTION_FLT_INEXACT_RESULT (STATUS_FLOAT_INEXACT_RESULT)
value EXCEPTION_FLT_INVALID_OPERATION (STATUS_FLOAT_INVALID_OPERATION)
value EXCEPTION_FLT_OVERFLOW (STATUS_FLOAT_OVERFLOW)
value EXCEPTION_FLT_STACK_CHECK (STATUS_FLOAT_STACK_CHECK)
value EXCEPTION_FLT_UNDERFLOW (STATUS_FLOAT_UNDERFLOW)
value EXCEPTION_GUARD_PAGE (STATUS_GUARD_PAGE_VIOLATION)
value EXCEPTION_ILLEGAL_INSTRUCTION (STATUS_ILLEGAL_INSTRUCTION)
value EXCEPTION_INT_DIVIDE_BY_ZERO (STATUS_INTEGER_DIVIDE_BY_ZERO)
value EXCEPTION_INT_OVERFLOW (STATUS_INTEGER_OVERFLOW)
value EXCEPTION_INVALID_DISPOSITION (STATUS_INVALID_DISPOSITION)
value EXCEPTION_INVALID_HANDLE (STATUS_INVALID_HANDLE)
value EXCEPTION_IN_PAGE_ERROR (STATUS_IN_PAGE_ERROR)
value EXCEPTION_MAXIMUM_PARAMETERS (15)
value EXCEPTION_NONCONTINUABLE_EXCEPTION (STATUS_NONCONTINUABLE_EXCEPTION)
value EXCEPTION_POSSIBLE_DEADLOCK (STATUS_POSSIBLE_DEADLOCK)
value EXCEPTION_PRIV_INSTRUCTION (STATUS_PRIVILEGED_INSTRUCTION)
value EXCEPTION_READ_FAULT (0)
value EXCEPTION_SINGLE_STEP (STATUS_SINGLE_STEP)
value EXCEPTION_STACK_OVERFLOW (STATUS_STACK_OVERFLOW)
value EXCEPTION_WRITE_FAULT (1)
value EXDEV (18)
value EXIT_FAILURE (1)
value EXIT_PROCESS_DEBUG_EVENT (5)
value EXIT_SUCCESS (0)
value EXIT_THREAD_DEBUG_EVENT (4)
value EXPENTRY (CALLBACK)
value EXTEND_IEPORT (2)
value EXTTEXTOUT (512)
value EXT_DEVICE_CAPS (4099)
value E_DRAW (VIEW_E_DRAW)
value FACILITY_AAF (18)
value FACILITY_ACCELERATOR (1536)
value FACILITY_ACS (20)
value FACILITY_ACTION_QUEUE (44)
value FACILITY_AUDCLNT (2185)
value FACILITY_AUDIO (102)
value FACILITY_AUDIOSTREAMING (1094)
value FACILITY_BACKGROUNDCOPY (32)
value FACILITY_BCD (57)
value FACILITY_BLB (120)
value FACILITY_BLBUI (128)
value FACILITY_BLB_CLI (121)
value FACILITY_BLUETOOTH_ATT (101)
value FACILITY_CERT (11)
value FACILITY_CMI (54)
value FACILITY_COMPLUS (17)
value FACILITY_CONFIGURATION (33)
value FACILITY_CONTROL (10)
value FACILITY_DAF (100)
value FACILITY_DEBUGGERS (176)
value FACILITY_DEFRAG (2304)
value FACILITY_DELIVERY_OPTIMIZATION (208)
value FACILITY_DEPLOYMENT_SERVICES_BINLSVC (261)
value FACILITY_DEPLOYMENT_SERVICES_CONTENT_PROVIDER (293)
value FACILITY_DEPLOYMENT_SERVICES_DRIVER_PROVISIONING (278)
value FACILITY_DEPLOYMENT_SERVICES_IMAGING (258)
value FACILITY_DEPLOYMENT_SERVICES_MANAGEMENT (259)
value FACILITY_DEPLOYMENT_SERVICES_MULTICAST_CLIENT (290)
value FACILITY_DEPLOYMENT_SERVICES_MULTICAST_SERVER (289)
value FACILITY_DEPLOYMENT_SERVICES_PXE (263)
value FACILITY_DEPLOYMENT_SERVICES_SERVER (257)
value FACILITY_DEPLOYMENT_SERVICES_TFTP (264)
value FACILITY_DEPLOYMENT_SERVICES_TRANSPORT_MANAGEMENT (272)
value FACILITY_DEPLOYMENT_SERVICES_UTIL (260)
value FACILITY_DEVICE_UPDATE_AGENT (135)
value FACILITY_DIRECTMUSIC (2168)
value FACILITY_DIRECTORYSERVICE (37)
value FACILITY_DISPATCH (2)
value FACILITY_DLS (153)
value FACILITY_DMSERVER (256)
value FACILITY_DPLAY (21)
value FACILITY_DRVSERVICING (136)
value FACILITY_DXCORE (2176)
value FACILITY_DXGI (2170)
value FACILITY_DXGI_DDI (2171)
value FACILITY_EAP (66)
value FACILITY_EAS (85)
value FACILITY_FVE (49)
value FACILITY_FWP (50)
value FACILITY_GAME (2340)
value FACILITY_GRAPHICS (38)
value FACILITY_HSP_SERVICES (296)
value FACILITY_HSP_SOFTWARE (297)
value FACILITY_HTTP (25)
value FACILITY_INPUT (64)
value FACILITY_INTERNET (12)
value FACILITY_IORING (70)
value FACILITY_ITF (4)
value FACILITY_JSCRIPT (2306)
value FACILITY_LEAP (2184)
value FACILITY_LINGUISTIC_SERVICES (305)
value FACILITY_MBN (84)
value FACILITY_MEDIASERVER (13)
value FACILITY_METADIRECTORY (35)
value FACILITY_MOBILE (1793)
value FACILITY_MSMQ (14)
value FACILITY_NAP (39)
value FACILITY_NDIS (52)
value FACILITY_NULL (0)
value FACILITY_OCP_UPDATE_AGENT (173)
value FACILITY_ONLINE_ID (134)
value FACILITY_OPC (81)
value FACILITY_PARSE (113)
value FACILITY_PIDGENX (2561)
value FACILITY_PIX (2748)
value FACILITY_PLA (48)
value FACILITY_POWERSHELL (84)
value FACILITY_PRESENTATION (2177)
value FACILITY_QUIC (65)
value FACILITY_RAS (83)
value FACILITY_RESTORE (256)
value FACILITY_RPC (1)
value FACILITY_SCARD (16)
value FACILITY_SCRIPT (112)
value FACILITY_SDIAG (60)
value FACILITY_SECURITY (9)
value FACILITY_SERVICE_FABRIC (1968)
value FACILITY_SETUPAPI (15)
value FACILITY_SHELL (39)
value FACILITY_SOS (160)
value FACILITY_SPP (256)
value FACILITY_SQLITE (1967)
value FACILITY_SSPI (9)
value FACILITY_STATEREPOSITORY (103)
value FACILITY_STATE_MANAGEMENT (34)
value FACILITY_STORAGE (3)
value FACILITY_SXS (23)
value FACILITY_SYNCENGINE (2050)
value FACILITY_TIERING (131)
value FACILITY_TPM_SERVICES (40)
value FACILITY_TPM_SOFTWARE (41)
value FACILITY_TTD (1490)
value FACILITY_UI (42)
value FACILITY_UMI (22)
value FACILITY_URT (19)
value FACILITY_USERMODE_COMMONLOG (26)
value FACILITY_USERMODE_FILTER_MANAGER (31)
value FACILITY_USERMODE_HNS (59)
value FACILITY_USERMODE_HYPERVISOR (53)
value FACILITY_USERMODE_LICENSING (234)
value FACILITY_USERMODE_SDBUS (2305)
value FACILITY_USERMODE_SPACES (231)
value FACILITY_USERMODE_VHD (58)
value FACILITY_USERMODE_VIRTUALIZATION (55)
value FACILITY_USERMODE_VOLMGR (56)
value FACILITY_USERMODE_VOLSNAP (130)
value FACILITY_USER_MODE_SECURITY_CORE (232)
value FACILITY_USN (129)
value FACILITY_UTC (1989)
value FACILITY_VISUALCPP (109)
value FACILITY_WEB (885)
value FACILITY_WEBSERVICES (61)
value FACILITY_WEB_SOCKET (886)
value FACILITY_WEP (2049)
value FACILITY_WER (27)
value FACILITY_WIA (33)
value FACILITY_WINCODEC_DWRITE_DWM (2200)
value FACILITY_WINDOWS (8)
value FACILITY_WINDOWSUPDATE (36)
value FACILITY_WINDOWS_CE (24)
value FACILITY_WINDOWS_DEFENDER (80)
value FACILITY_WINDOWS_SETUP (48)
value FACILITY_WINDOWS_STORE (63)
value FACILITY_WINML (2192)
value FACILITY_WINPE (61)
value FACILITY_WINRM (51)
value FACILITY_WMAAECMA (1996)
value FACILITY_WPN (62)
value FACILITY_WSBAPP (122)
value FACILITY_WSB_ONLINE (133)
value FACILITY_XAML (43)
value FACILITY_XBOX (2339)
value FACILITY_XPS (82)
value FALSE (0)
value FAPPCOMMAND_KEY (0)
value FAST_FAIL_ADMINLESS_ACCESS_DENIED (55)
value FAST_FAIL_APCS_DISABLED (32)
value FAST_FAIL_CAST_GUARD (65)
value FAST_FAIL_CERTIFICATION_FAILURE (20)
value FAST_FAIL_CONTROL_INVALID_RETURN_ADDRESS (57)
value FAST_FAIL_CORRUPT_LIST_ENTRY (3)
value FAST_FAIL_CRYPTO_LIBRARY (22)
value FAST_FAIL_DEPRECATED_SERVICE_INVOKED (27)
value FAST_FAIL_DLOAD_PROTECTION_FAILURE (25)
value FAST_FAIL_ENCLAVE_CALL_FAILURE (53)
value FAST_FAIL_ETW_CORRUPTION (61)
value FAST_FAIL_FATAL_APP_EXIT (7)
value FAST_FAIL_FLAGS_CORRUPTION (59)
value FAST_FAIL_GS_COOKIE_INIT (6)
value FAST_FAIL_GUARD_EXPORT_SUPPRESSION_FAILURE (46)
value FAST_FAIL_GUARD_ICALL_CHECK_FAILURE (10)
value FAST_FAIL_GUARD_ICALL_CHECK_FAILURE_XFG (64)
value FAST_FAIL_GUARD_ICALL_CHECK_SUPPRESSED (31)
value FAST_FAIL_GUARD_JUMPTABLE (37)
value FAST_FAIL_GUARD_SS_FAILURE (44)
value FAST_FAIL_GUARD_WRITE_CHECK_FAILURE (11)
value FAST_FAIL_HEAP_METADATA_CORRUPTION (50)
value FAST_FAIL_HOST_VISIBILITY_CHANGE (66)
value FAST_FAIL_INCORRECT_STACK (4)
value FAST_FAIL_INVALID_ARG (5)
value FAST_FAIL_INVALID_BALANCED_TREE (29)
value FAST_FAIL_INVALID_BUFFER_ACCESS (28)
value FAST_FAIL_INVALID_CALL_IN_DLL_CALLOUT (23)
value FAST_FAIL_INVALID_CONTROL_STACK (47)
value FAST_FAIL_INVALID_DISPATCH_CONTEXT (39)
value FAST_FAIL_INVALID_EXCEPTION_CHAIN (21)
value FAST_FAIL_INVALID_FIBER_SWITCH (12)
value FAST_FAIL_INVALID_FILE_OPERATION (42)
value FAST_FAIL_INVALID_FLS_DATA (70)
value FAST_FAIL_INVALID_IAT (49)
value FAST_FAIL_INVALID_IDLE_STATE (33)
value FAST_FAIL_INVALID_IMAGE_BASE (24)
value FAST_FAIL_INVALID_JUMP_BUFFER (18)
value FAST_FAIL_INVALID_LOCK_STATE (36)
value FAST_FAIL_INVALID_LONGJUMP_TARGET (38)
value FAST_FAIL_INVALID_NEXT_THREAD (30)
value FAST_FAIL_INVALID_PFN (63)
value FAST_FAIL_INVALID_REFERENCE_COUNT (14)
value FAST_FAIL_INVALID_SET_OF_CONTEXT (13)
value FAST_FAIL_INVALID_SYSCALL_NUMBER (41)
value FAST_FAIL_INVALID_THREAD (40)
value FAST_FAIL_KERNEL_CET_SHADOW_STACK_ASSIST (67)
value FAST_FAIL_LEGACY_GS_VIOLATION (0)
value FAST_FAIL_LOADER_CONTINUITY_FAILURE (45)
value FAST_FAIL_LOW_LABEL_ACCESS_DENIED (52)
value FAST_FAIL_LPAC_ACCESS_DENIED (43)
value FAST_FAIL_MRDATA_MODIFIED (19)
value FAST_FAIL_MRDATA_PROTECTION_FAILURE (34)
value FAST_FAIL_NTDLL_PATCH_FAILED (69)
value FAST_FAIL_PATCH_CALLBACK_FAILED (68)
value FAST_FAIL_PAYLOAD_RESTRICTION_VIOLATION (51)
value FAST_FAIL_RANGE_CHECK_FAILURE (8)
value FAST_FAIL_RIO_ABORT (62)
value FAST_FAIL_SET_CONTEXT_DENIED (48)
value FAST_FAIL_STACK_COOKIE_CHECK_FAILURE (2)
value FAST_FAIL_UNEXPECTED_CALL (56)
value FAST_FAIL_UNEXPECTED_HEAP_EXCEPTION (35)
value FAST_FAIL_UNEXPECTED_HOST_BEHAVIOR (58)
value FAST_FAIL_UNHANDLED_LSS_EXCEPTON (54)
value FAST_FAIL_UNSAFE_EXTENSION_CALL (26)
value FAST_FAIL_UNSAFE_REGISTRY_ACCESS (9)
value FAST_FAIL_VEH_CORRUPTION (60)
value FAST_FAIL_VTGUARD_CHECK_FAILURE (1)
value FD_ACCEPT_BIT (3)
value FD_ADDRESS_LIST_CHANGE_BIT (9)
value FD_CLOSE_BIT (5)
value FD_CONNECT_BIT (4)
value FD_GROUP_QOS_BIT (7)
value FD_MAX_EVENTS (10)
value FD_OOB_BIT (2)
value FD_QOS_BIT (6)
value FD_READ_BIT (0)
value FD_ROUTING_INTERFACE_CHANGE_BIT (8)
value FD_SETSIZE (64)
value FD_WRITE_BIT (1)
value FEATURESETTING_CUSTPAPER (3)
value FEATURESETTING_MIRROR (4)
value FEATURESETTING_NEGATIVE (5)
value FEATURESETTING_NUP (0)
value FEATURESETTING_OUTPUT (1)
value FEATURESETTING_PROTOCOL (6)
value FEATURESETTING_PSLEVEL (2)
value FILENAME_MAX (260)
value FILEOKSTRING (FILEOKSTRINGA)
value FILEOPENORD (1536)
value FILESYSTEM_STATISTICS_TYPE_EXFAT (3)
value FILESYSTEM_STATISTICS_TYPE_FAT (2)
value FILESYSTEM_STATISTICS_TYPE_NTFS (1)
value FILESYSTEM_STATISTICS_TYPE_REFS (4)
value FILE_ANY_ACCESS (0)
value FILE_BEGIN (0)
value FILE_CURRENT (1)
value FILE_DIR_DISALLOWED (9)
value FILE_ENCRYPTABLE (0)
value FILE_END (2)
value FILE_IS_ENCRYPTED (1)
value FILE_MAP_ALL_ACCESS (SECTION_ALL_ACCESS)
value FILE_MAP_EXECUTE (SECTION_MAP_EXECUTE_EXPLICIT)
value FILE_MAP_READ (SECTION_MAP_READ)
value FILE_MAP_WRITE (SECTION_MAP_WRITE)
value FILE_NAME_FLAG_HARDLINK (0)
value FILE_READ_ONLY (8)
value FILE_ROOT_DIR (3)
value FILE_SYSTEM_ATTR (2)
value FILE_SYSTEM_DIR (4)
value FILE_SYSTEM_NOT_SUPPORT (6)
value FILE_UNKNOWN (5)
value FILE_USER_DISALLOWED (7)
value FINDDLGORD (1540)
value FINDMSGSTRING (FINDMSGSTRINGA)
value FIXED_PITCH (1)
value FLASHW_STOP (0)
value FLOODFILLBORDER (0)
value FLOODFILLSURFACE (1)
value FLS_MAXIMUM_AVAILABLE (4080)
value FLUSHOUTPUT (6)
value FMTID_NULL (GUID_NULL)
value FONTDLGORD (1542)
value FONTMAPPER_MAX (10)
value FOPEN_MAX (20)
value FRAME_FPO (0)
value FRAME_NONFPO (3)
value FRAME_TRAP (1)
value FRAME_TSS (2)
value FRS_ERR_AUTHENTICATION (8008L)
value FRS_ERR_CHILD_TO_PARENT_COMM (8011L)
value FRS_ERR_INSUFFICIENT_PRIV (8007L)
value FRS_ERR_INTERNAL (8005L)
value FRS_ERR_INTERNAL_API (8004L)
value FRS_ERR_INVALID_API_SEQUENCE (8001L)
value FRS_ERR_INVALID_SERVICE_PARAMETER (8017L)
value FRS_ERR_PARENT_AUTHENTICATION (8010L)
value FRS_ERR_PARENT_INSUFFICIENT_PRIV (8009L)
value FRS_ERR_PARENT_TO_CHILD_COMM (8012L)
value FRS_ERR_SERVICE_COMM (8006L)
value FRS_ERR_STARTING_SERVICE (8002L)
value FRS_ERR_STOPPING_SERVICE (8003L)
value FRS_ERR_SYSVOL_DEMOTE (8016L)
value FRS_ERR_SYSVOL_IS_BUSY (8015L)
value FRS_ERR_SYSVOL_POPULATE (8013L)
value FRS_ERR_SYSVOL_POPULATE_TIMEOUT (8014L)
value FSCTL_MARK_AS_SYSTEM_HIVE (FSCTL_SET_BOOTLOADER_ACCESSED)
value FS_CASE_IS_PRESERVED (FILE_CASE_PRESERVED_NAMES)
value FS_CASE_SENSITIVE (FILE_CASE_SENSITIVE_SEARCH)
value FS_FILE_COMPRESSION (FILE_FILE_COMPRESSION)
value FS_FILE_ENCRYPTION (FILE_SUPPORTS_ENCRYPTION)
value FS_PERSISTENT_ACLS (FILE_PERSISTENT_ACLS)
value FS_UNICODE_STORED_ON_DISK (FILE_UNICODE_ON_DISK)
value FS_VOL_IS_COMPRESSED (FILE_VOLUME_IS_COMPRESSED)
value FVIRTKEY (TRUE)
value FW_BLACK (FW_HEAVY)
value FW_BOLD (700)
value FW_DEMIBOLD (FW_SEMIBOLD)
value FW_DONTCARE (0)
value FW_EXTRABOLD (800)
value FW_EXTRALIGHT (200)
value FW_HEAVY (900)
value FW_LIGHT (300)
value FW_MEDIUM (500)
value FW_NORMAL (400)
value FW_REGULAR (FW_NORMAL)
value FW_SEMIBOLD (600)
value FW_THIN (100)
value FW_ULTRABOLD (FW_EXTRABOLD)
value FW_ULTRALIGHT (FW_EXTRALIGHT)
value GA_PARENT (1)
value GA_ROOT (2)
value GA_ROOTOWNER (3)
value GCPCLASS_ARABIC (2)
value GCPCLASS_HEBREW (2)
value GCPCLASS_LATIN (1)
value GCPCLASS_LATINNUMBER (5)
value GCPCLASS_LATINNUMERICSEPARATOR (7)
value GCPCLASS_LATINNUMERICTERMINATOR (6)
value GCPCLASS_LOCALNUMBER (4)
value GCPCLASS_NEUTRAL (3)
value GCPCLASS_NUMERICSEPARATOR (8)
value GC_ROLLOVER (GC_PRESSANDTAP)
value GDIPLUS_TS_QUERYVER (4122)
value GDIPLUS_TS_RECORD (4123)
value GDI_MAX_OBJ_TYPE (GDI_OBJ_LAST)
value GDI_MIN_OBJ_TYPE (OBJ_PEN)
value GDI_OBJ_LAST (OBJ_COLORSPACE)
value GEO_NAME_USER_DEFAULT (NULL)
value GESTURECONFIGMAXCOUNT (256)
value GETCOLORTABLE (5)
value GETDEVICEUNITS (42)
value GETEXTENDEDTEXTMETRICS (256)
value GETEXTENTTABLE (257)
value GETFACENAME (513)
value GETPAIRKERNTABLE (258)
value GETPENWIDTH (16)
value GETPHYSPAGESIZE (12)
value GETPRINTINGOFFSET (13)
value GETSCALINGFACTOR (14)
value GETSETPAPERBINS (29)
value GETSETPAPERMETRICS (35)
value GETSETPRINTORIENT (30)
value GETSETSCREENPARAMS (3072)
value GETTECHNOLGY (20)
value GETTECHNOLOGY (20)
value GETTRACKKERNTABLE (259)
value GETVECTORBRUSHSIZE (27)
value GETVECTORPENSIZE (26)
value GET_MOUSEORKEY_LPARAM (GET_DEVICE_LPARAM)
value GET_PS_FEATURESETTING (4121)
value GET_TAPE_DRIVE_INFORMATION (1)
value GET_TAPE_MEDIA_INFORMATION (0)
value GGI_MARK_NONEXISTING_GLYPHS (0cX0001)
value GGO_BEZIER (3)
value GGO_BITMAP (1)
value GGO_METRICS (0)
value GGO_NATIVE (2)
value GIDC_ARRIVAL (1)
value GIDC_REMOVAL (2)
value GID_BEGIN (1)
value GID_END (2)
value GID_PAN (4)
value GID_PRESSANDTAP (7)
value GID_ROLLOVER (GID_PRESSANDTAP)
value GID_ROTATE (5)
value GID_TWOFINGERTAP (6)
value GID_ZOOM (3)
value GMEM_LOWER (GMEM_NOT_BANKED)
value GMMP_USE_DISPLAY_POINTS (1)
value GMMP_USE_HIGH_RESOLUTION_POINTS (2)
value GM_ADVANCED (2)
value GM_COMPATIBLE (1)
value GM_LAST (2)
value GRAY_BRUSH (2)
value GREEK_CHARSET (161)
value GR_GDIOBJECTS (0)
value GR_GDIOBJECTS_PEAK (2)
value GR_USEROBJECTS (1)
value GR_USEROBJECTS_PEAK (4)
value GUID_CLASS_COMPORT (GUID_DEVINTERFACE_COMPORT)
value GUID_SERENUM_BUS_ENUMERATOR (GUID_DEVINTERFACE_SERENUM_BUS_ENUMERATOR)
value GW_CHILD (5)
value GW_ENABLEDPOPUP (6)
value GW_HWNDFIRST (0)
value GW_HWNDLAST (1)
value GW_HWNDNEXT (2)
value GW_HWNDPREV (3)
value GW_MAX (6)
value GW_OWNER (4)
value HALFTONE (4)
value HANGEUL_CHARSET (129)
value HANGUL_CHARSET (129)
value HCBT_ACTIVATE (5)
value HCBT_CLICKSKIPPED (6)
value HCBT_CREATEWND (3)
value HCBT_DESTROYWND (4)
value HCBT_KEYSKIPPED (7)
value HCBT_MINMAX (1)
value HCBT_MOVESIZE (0)
value HCBT_QS (2)
value HCBT_SETFOCUS (9)
value HCBT_SYSCOMMAND (8)
value HC_ACTION (0)
value HC_GETNEXT (1)
value HC_NOREM (HC_NOREMOVE)
value HC_NOREMOVE (3)
value HC_SKIP (2)
value HC_SYSMODALOFF (5)
value HC_SYSMODALON (4)
value HEAP_OPTIMIZE_RESOURCES_CURRENT_VERSION (1)
value HEAP_TAG_SHIFT (18)
value HEBREW_CHARSET (177)
value HELPMSGSTRING (HELPMSGSTRINGA)
value HIDE_WINDOW (0)
value HIGH_LEVEL (15)
value HINSTANCE_ERROR (32)
value HIST_NO_OF_BUCKETS (24)
value HKL_NEXT (1)
value HKL_PREV (0)
value HOLLOW_BRUSH (NULL_BRUSH)
value HORZRES (8)
value HORZSIZE (4)
value HOST_NOT_FOUND (WSAHOST_NOT_FOUND)
value HSHELL_ACCESSIBILITYSTATE (11)
value HSHELL_ACTIVATESHELLWINDOW (3)
value HSHELL_APPCOMMAND (12)
value HSHELL_ENDTASK (10)
value HSHELL_GETMINRECT (5)
value HSHELL_LANGUAGE (8)
value HSHELL_MONITORCHANGED (16)
value HSHELL_REDRAW (6)
value HSHELL_SYSMENU (9)
value HSHELL_TASKMAN (7)
value HSHELL_WINDOWACTIVATED (4)
value HSHELL_WINDOWCREATED (1)
value HSHELL_WINDOWDESTROYED (2)
value HSHELL_WINDOWREPLACED (13)
value HSHELL_WINDOWREPLACING (14)
value HS_API_MAX (12)
value HS_BDIAGONAL (3)
value HS_CROSS (4)
value HS_DIAGCROSS (5)
value HS_FDIAGONAL (2)
value HS_HORIZONTAL (0)
value HS_VERTICAL (1)
value HTBORDER (18)
value HTBOTTOM (15)
value HTBOTTOMLEFT (16)
value HTBOTTOMRIGHT (17)
value HTCAPTION (2)
value HTCLIENT (1)
value HTCLOSE (20)
value HTGROWBOX (4)
value HTHELP (21)
value HTHSCROLL (6)
value HTLEFT (10)
value HTMAXBUTTON (9)
value HTMENU (5)
value HTMINBUTTON (8)
value HTNOWHERE (0)
value HTOBJECT (19)
value HTREDUCE (HTMINBUTTON)
value HTRIGHT (11)
value HTSIZE (HTGROWBOX)
value HTSIZEFIRST (HTLEFT)
value HTSIZELAST (HTBOTTOMRIGHT)
value HTSYSMENU (3)
value HTTOP (12)
value HTTOPLEFT (13)
value HTTOPRIGHT (14)
value HTVSCROLL (7)
value HTZOOM (HTMAXBUTTON)
value HW_PROFILE_GUIDLEN (39)
value ICMENUMPROC (ICMENUMPROCA)
value ICM_ADDPROFILE (1)
value ICM_DELETEPROFILE (2)
value ICM_DONE_OUTSIDEDC (4)
value ICM_OFF (1)
value ICM_ON (2)
value ICM_QUERY (3)
value ICM_QUERYMATCH (7)
value ICM_QUERYPROFILE (3)
value ICM_REGISTERICMATCHER (5)
value ICM_SETDEFAULTPROFILE (4)
value ICM_UNREGISTERICMATCHER (6)
value ICON_BIG (1)
value ICON_SMALL (0)
value IDABORT (3)
value IDANI_CAPTION (3)
value IDANI_OPEN (1)
value IDCANCEL (2)
value IDCLOSE (8)
value IDCONTINUE (11)
value IDC_MANAGE_LINK (1592)
value IDENTIFY_BUFFER_SIZE (512)
value IDHELP (9)
value IDH_CANCEL (28444)
value IDH_GENERIC_HELP_BUTTON (28442)
value IDH_HELP (28445)
value IDH_MISSING_CONTEXT (28441)
value IDH_NO_HELP (28440)
value IDH_OK (28443)
value IDIGNORE (5)
value IDI_ERROR (IDI_HAND)
value IDI_INFORMATION (IDI_ASTERISK)
value IDI_WARNING (IDI_EXCLAMATION)
value IDNO (7)
value IDOK (1)
value IDRETRY (4)
value IDTIMEOUT (32000)
value IDTRYAGAIN (10)
value IDYES (6)
value IFX_RSA_KEYGEN_VUL_NOT_AFFECTED (0)
value IGNORE (0)
value IID_NULL (GUID_NULL)
value ILLUMINANT_A (1)
value ILLUMINANT_B (2)
value ILLUMINANT_C (3)
value ILLUMINANT_DAYLIGHT (ILLUMINANT_C)
value ILLUMINANT_DEVICE_DEFAULT (0)
value ILLUMINANT_FLUORESCENT (ILLUMINANT_F2)
value ILLUMINANT_MAX_INDEX (ILLUMINANT_F2)
value ILLUMINANT_NTSC (ILLUMINANT_C)
value ILLUMINANT_TUNGSTEN (ILLUMINANT_A)
value IMAGE_ARCHIVE_START_SIZE (8)
value IMAGE_BITMAP (0)
value IMAGE_COMDAT_SELECT_ANY (2)
value IMAGE_COMDAT_SELECT_ASSOCIATIVE (5)
value IMAGE_COMDAT_SELECT_EXACT_MATCH (4)
value IMAGE_COMDAT_SELECT_LARGEST (6)
value IMAGE_COMDAT_SELECT_NEWEST (7)
value IMAGE_COMDAT_SELECT_NODUPLICATES (1)
value IMAGE_COMDAT_SELECT_SAME_SIZE (3)
value IMAGE_CURSOR (2)
value IMAGE_DEBUG_MISC_EXENAME (1)
value IMAGE_DEBUG_TYPE_BBT (IMAGE_DEBUG_TYPE_RESERVED10)
value IMAGE_DEBUG_TYPE_BORLAND (9)
value IMAGE_DEBUG_TYPE_CLSID (11)
value IMAGE_DEBUG_TYPE_CODEVIEW (2)
value IMAGE_DEBUG_TYPE_COFF (1)
value IMAGE_DEBUG_TYPE_EXCEPTION (5)
value IMAGE_DEBUG_TYPE_EX_DLLCHARACTERISTICS (20)
value IMAGE_DEBUG_TYPE_FIXUP (6)
value IMAGE_DEBUG_TYPE_FPO (3)
value IMAGE_DEBUG_TYPE_ILTCG (14)
value IMAGE_DEBUG_TYPE_MISC (4)
value IMAGE_DEBUG_TYPE_MPX (15)
value IMAGE_DEBUG_TYPE_OMAP_FROM_SRC (8)
value IMAGE_DEBUG_TYPE_OMAP_TO_SRC (7)
value IMAGE_DEBUG_TYPE_POGO (13)
value IMAGE_DEBUG_TYPE_REPRO (16)
value IMAGE_DEBUG_TYPE_SPGO (18)
value IMAGE_DEBUG_TYPE_UNKNOWN (0)
value IMAGE_DEBUG_TYPE_VC_FEATURE (12)
value IMAGE_DIRECTORY_ENTRY_ARCHITECTURE (7)
value IMAGE_DIRECTORY_ENTRY_BASERELOC (5)
value IMAGE_DIRECTORY_ENTRY_BOUND_IMPORT (11)
value IMAGE_DIRECTORY_ENTRY_COM_DESCRIPTOR (14)
value IMAGE_DIRECTORY_ENTRY_DEBUG (6)
value IMAGE_DIRECTORY_ENTRY_DELAY_IMPORT (13)
value IMAGE_DIRECTORY_ENTRY_EXCEPTION (3)
value IMAGE_DIRECTORY_ENTRY_EXPORT (0)
value IMAGE_DIRECTORY_ENTRY_GLOBALPTR (8)
value IMAGE_DIRECTORY_ENTRY_IAT (12)
value IMAGE_DIRECTORY_ENTRY_IMPORT (1)
value IMAGE_DIRECTORY_ENTRY_LOAD_CONFIG (10)
value IMAGE_DIRECTORY_ENTRY_RESOURCE (2)
value IMAGE_DIRECTORY_ENTRY_SECURITY (4)
value IMAGE_DIRECTORY_ENTRY_TLS (9)
value IMAGE_ENCLAVE_LONG_ID_LENGTH (ENCLAVE_LONG_ID_LENGTH)
value IMAGE_ENCLAVE_SHORT_ID_LENGTH (ENCLAVE_SHORT_ID_LENGTH)
value IMAGE_ENHMETAFILE (3)
value IMAGE_FILE_MACHINE_UNKNOWN (0)
value IMAGE_FUNCTION_OVERRIDE_INVALID (0)
value IMAGE_GUARD_CF_FUNCTION_TABLE_SIZE_SHIFT (28)
value IMAGE_ICON (1)
value IMAGE_NT_OPTIONAL_HDR_MAGIC (IMAGE_NT_OPTIONAL_HDR64_MAGIC)
value IMAGE_NUMBEROF_DIRECTORY_ENTRIES (16)
value IMAGE_ORDINAL_FLAG (IMAGE_ORDINAL_FLAG64)
value IMAGE_POLICY_METADATA_VERSION (1)
value IMAGE_REL_BASED_ABSOLUTE (0)
value IMAGE_REL_BASED_HIGH (1)
value IMAGE_REL_BASED_HIGHADJ (4)
value IMAGE_REL_BASED_HIGHLOW (3)
value IMAGE_REL_BASED_LOW (2)
value IMAGE_REL_BASED_MIPS_JMPADDR (5)
value IMAGE_REL_BASED_RESERVED (6)
value IMAGE_SIZEOF_ARCHIVE_MEMBER_HDR (60)
value IMAGE_SIZEOF_FILE_HEADER (20)
value IMAGE_SIZEOF_SECTION_HEADER (40)
value IMAGE_SIZEOF_SHORT_NAME (8)
value IMAGE_SIZEOF_SYMBOL (18)
value IMAGE_SUBSYSTEM_EFI_APPLICATION (10)
value IMAGE_SUBSYSTEM_EFI_BOOT_SERVICE_DRIVER (11)
value IMAGE_SUBSYSTEM_EFI_ROM (13)
value IMAGE_SUBSYSTEM_EFI_RUNTIME_DRIVER (12)
value IMAGE_SUBSYSTEM_NATIVE (1)
value IMAGE_SUBSYSTEM_NATIVE_WINDOWS (8)
value IMAGE_SUBSYSTEM_POSIX_CUI (7)
value IMAGE_SUBSYSTEM_UNKNOWN (0)
value IMAGE_SUBSYSTEM_WINDOWS_BOOT_APPLICATION (16)
value IMAGE_SUBSYSTEM_WINDOWS_CE_GUI (9)
value IMAGE_SUBSYSTEM_WINDOWS_CUI (3)
value IMAGE_SUBSYSTEM_WINDOWS_GUI (2)
value IMAGE_SUBSYSTEM_XBOX (14)
value IMAGE_SUBSYSTEM_XBOX_CODE_CATALOG (17)
value IMAGE_SYM_DTYPE_ARRAY (3)
value IMAGE_SYM_DTYPE_FUNCTION (2)
value IMAGE_SYM_DTYPE_NULL (0)
value IMAGE_SYM_DTYPE_POINTER (1)
value IMAGE_SYM_SECTION_MAX_EX (MAXLONG)
value IMAGE_WEAK_EXTERN_ANTI_DEPENDENCY (4)
value IMAGE_WEAK_EXTERN_SEARCH_ALIAS (3)
value IMAGE_WEAK_EXTERN_SEARCH_LIBRARY (2)
value IMAGE_WEAK_EXTERN_SEARCH_NOLIBRARY (1)
value IMEMENUITEM_STRING_SIZE (80)
value IME_CMODE_CHINESE (IME_CMODE_NATIVE)
value IME_CMODE_HANGEUL (IME_CMODE_NATIVE)
value IME_CMODE_HANGUL (IME_CMODE_NATIVE)
value IME_CMODE_JAPANESE (IME_CMODE_NATIVE)
value IME_CONFIG_GENERAL (1)
value IME_CONFIG_REGISTERWORD (2)
value IME_CONFIG_SELECTDICTIONARY (3)
value IMFS_CHECKED (MFS_CHECKED)
value IMFS_DEFAULT (MFS_DEFAULT)
value IMFS_DISABLED (MFS_DISABLED)
value IMFS_ENABLED (MFS_ENABLED)
value IMFS_GRAYED (MFS_GRAYED)
value IMFS_HILITE (MFS_HILITE)
value IMFS_UNCHECKED (MFS_UNCHECKED)
value IMFS_UNHILITE (MFS_UNHILITE)
value IMPLINK_HIGHEXPER (158)
value IMPLINK_IP (155)
value IMPLINK_LOWEXPER (156)
value INCL_WINSOCK_API_PROTOTYPES (1)
value INCL_WINSOCK_API_TYPEDEFS (0)
value INDEXID_CONTAINER (0)
value INDEXID_OBJECT (0)
value INET_E_DEFAULT_ACTION (INET_E_USE_DEFAULT_PROTOCOLHANDLER)
value INET_E_ERROR_LAST (INET_E_DOWNLOAD_BLOCKED_BY_CSP)
value INIT_ONCE_ASYNC (RTL_RUN_ONCE_ASYNC)
value INIT_ONCE_CHECK_ONLY (RTL_RUN_ONCE_CHECK_ONLY)
value INIT_ONCE_CTX_RESERVED_BITS (RTL_RUN_ONCE_CTX_RESERVED_BITS)
value INIT_ONCE_INIT_FAILED (RTL_RUN_ONCE_INIT_FAILED)
value INIT_ONCE_STATIC_INIT (RTL_RUN_ONCE_INIT)
value INPUT_HARDWARE (2)
value INPUT_KEYBOARD (1)
value INPUT_MOUSE (0)
value INT_MAX (2147483647)
value IN_CLASSA_MAX (128)
value IN_CLASSA_NSHIFT (24)
value IN_CLASSB_MAX (65536)
value IN_CLASSB_NSHIFT (16)
value IN_CLASSC_NSHIFT (8)
value IN_CLASSD_NSHIFT (28)
value IOCTL_CHANGER_BASE (FILE_DEVICE_CHANGER)
value IOCTL_DISK_BASE (FILE_DEVICE_DISK)
value IOCTL_SCMBUS_BASE (FILE_DEVICE_PERSISTENT_MEMORY)
value IOCTL_STORAGE_BASE (FILE_DEVICE_MASS_STORAGE)
value IOCTL_STORAGE_BC_VERSION (1)
value IO_QOS_MAX_RESERVATION (1000000000ULL)
value IO_REPARSE_TAG_RESERVED_RANGE (IO_REPARSE_TAG_RESERVED_TWO)
value IPPORT_BIFFUDP (512)
value IPPORT_CHARGEN (19)
value IPPORT_CMDSERVER (514)
value IPPORT_DAYTIME (13)
value IPPORT_DISCARD (9)
value IPPORT_ECHO (7)
value IPPORT_EFSSERVER (520)
value IPPORT_EPMAP (135)
value IPPORT_EXECSERVER (512)
value IPPORT_FINGER (79)
value IPPORT_FTP (21)
value IPPORT_FTP_DATA (20)
value IPPORT_HTTPS (443)
value IPPORT_IMAP (143)
value IPPORT_LDAP (389)
value IPPORT_LOGINSERVER (513)
value IPPORT_MICROSOFT_DS (445)
value IPPORT_MSP (18)
value IPPORT_MTP (57)
value IPPORT_NAMESERVER (42)
value IPPORT_NETBIOS_DGM (138)
value IPPORT_NETBIOS_NS (137)
value IPPORT_NETBIOS_SSN (139)
value IPPORT_NETSTAT (15)
value IPPORT_NTP (123)
value IPPORT_QOTD (17)
value IPPORT_REGISTERED_MIN (IPPORT_RESERVED)
value IPPORT_RESERVED (1024)
value IPPORT_RJE (77)
value IPPORT_ROUTESERVER (520)
value IPPORT_SMTP (25)
value IPPORT_SNMP (161)
value IPPORT_SNMP_TRAP (162)
value IPPORT_SUPDUP (95)
value IPPORT_SYSTAT (11)
value IPPORT_TCPMUX (1)
value IPPORT_TELNET (23)
value IPPORT_TFTP (69)
value IPPORT_TIMESERVER (37)
value IPPORT_TTYLINK (87)
value IPPORT_WHOIS (43)
value IPPORT_WHOSERVER (513)
value IPPROTO_IP (0)
value JOB_CONTROL_CANCEL (3)
value JOB_CONTROL_DELETE (5)
value JOB_CONTROL_LAST_PAGE_EJECTED (7)
value JOB_CONTROL_PAUSE (1)
value JOB_CONTROL_RELEASE (9)
value JOB_CONTROL_RESTART (4)
value JOB_CONTROL_RESUME (2)
value JOB_CONTROL_RETAIN (8)
value JOB_CONTROL_SEND_TOAST (10)
value JOB_CONTROL_SENT_TO_PRINTER (6)
value JOB_OBJECT_LIMIT_CPU_RATE_CONTROL (JOB_OBJECT_LIMIT_RATE_CONTROL)
value JOB_OBJECT_LIMIT_JOB_MEMORY_HIGH (JOB_OBJECT_LIMIT_JOB_MEMORY)
value JOB_OBJECT_MSG_ABNORMAL_EXIT_PROCESS (8)
value JOB_OBJECT_MSG_ACTIVE_PROCESS_LIMIT (3)
value JOB_OBJECT_MSG_ACTIVE_PROCESS_ZERO (4)
value JOB_OBJECT_MSG_END_OF_JOB_TIME (1)
value JOB_OBJECT_MSG_END_OF_PROCESS_TIME (2)
value JOB_OBJECT_MSG_EXIT_PROCESS (7)
value JOB_OBJECT_MSG_JOB_CYCLE_TIME_LIMIT (12)
value JOB_OBJECT_MSG_JOB_MEMORY_LIMIT (10)
value JOB_OBJECT_MSG_MAXIMUM (13)
value JOB_OBJECT_MSG_MINIMUM (1)
value JOB_OBJECT_MSG_NEW_PROCESS (6)
value JOB_OBJECT_MSG_NOTIFICATION_LIMIT (11)
value JOB_OBJECT_MSG_PROCESS_MEMORY_LIMIT (9)
value JOB_OBJECT_MSG_SILO_TERMINATED (13)
value JOB_OBJECT_NET_RATE_CONTROL_MAX_DSCP_TAG (64)
value JOB_OBJECT_POST_AT_END_OF_JOB (1)
value JOB_OBJECT_TERMINATE_AT_END_OF_JOB (0)
value JOB_POSITION_UNSPECIFIED (0)
value JOHAB_CHARSET (130)
value JOYERR_BASE (160)
value JOY_POVBACKWARD (18000)
value JOY_POVFORWARD (0)
value JOY_POVLEFT (27000)
value JOY_POVRIGHT (9000)
value KL_NAMELENGTH (9)
value KP_ADMIN_PIN (31)
value KP_ALGID (7)
value KP_BLOCKLEN (8)
value KP_CERTIFICATE (26)
value KP_CLEAR_KEY (27)
value KP_CLIENT_RANDOM (21)
value KP_CMS_DH_KEY_INFO (38)
value KP_CMS_KEY_INFO (37)
value KP_EFFECTIVE_KEYLEN (19)
value KP_G (12)
value KP_GET_USE_COUNT (42)
value KP_HIGHEST_VERSION (41)
value KP_INFO (18)
value KP_IV (1)
value KP_KEYEXCHANGE_PIN (32)
value KP_KEYLEN (9)
value KP_KEYVAL (30)
value KP_MODE (4)
value KP_MODE_BITS (5)
value KP_OAEP_PARAMS (36)
value KP_P (11)
value KP_PADDING (3)
value KP_PERMISSIONS (6)
value KP_PIN_ID (43)
value KP_PIN_INFO (44)
value KP_PRECOMP_SHA (25)
value KP_PREHASH (34)
value KP_PUB_EX_LEN (28)
value KP_PUB_EX_VAL (29)
value KP_PUB_PARAMS (39)
value KP_Q (13)
value KP_RA (16)
value KP_RB (17)
value KP_ROUNDS (35)
value KP_RP (23)
value KP_SALT (2)
value KP_SALT_EX (10)
value KP_SCHANNEL_ALG (20)
value KP_SERVER_RANDOM (22)
value KP_SIGNATURE_PIN (33)
value KP_VERIFY_PARAMS (40)
value KP_X (14)
value KP_Y (15)
value KTM_MARSHAL_BLOB_VERSION_MAJOR (1)
value KTM_MARSHAL_BLOB_VERSION_MINOR (1)
value LANGGROUPLOCALE_ENUMPROC (LANGGROUPLOCALE_ENUMPROCA)
value LANGUAGEGROUP_ENUMPROC (LANGUAGEGROUP_ENUMPROCA)
value LAYERED_PROTOCOL (0)
value LBN_DBLCLK (2)
value LBN_KILLFOCUS (5)
value LBN_SELCANCEL (3)
value LBN_SELCHANGE (1)
value LBN_SETFOCUS (4)
value LBSELCHSTRING (LBSELCHSTRINGA)
value LB_CTLCODE (0cL)
value LB_OKAY (0)
value LC_INTERIORS (128)
value LC_MARKER (4)
value LC_NONE (0)
value LC_POLYLINE (2)
value LC_POLYMARKER (8)
value LC_STYLED (32)
value LC_WIDE (16)
value LC_WIDESTYLED (64)
value LF_FACESIZE (32)
value LF_FULLFACESIZE (64)
value LINECAPS (30)
value LOAD_DLL_DEBUG_EVENT (6)
value LOCALE_ALL (0)
value LOCALE_ENUMPROC (LOCALE_ENUMPROCA)
value LOCALE_ICOUNTRY (LOCALE_IDIALINGCODE)
value LOCALE_NAME_MAX_LENGTH (85)
value LOCALE_NAME_USER_DEFAULT (NULL)
value LOCALE_SCOUNTRY (LOCALE_SLOCALIZEDCOUNTRYNAME)
value LOCALE_SENGCOUNTRY (LOCALE_SENGLISHCOUNTRYNAME)
value LOCALE_SENGLANGUAGE (LOCALE_SENGLISHLANGUAGENAME)
value LOCALE_SLANGDISPLAYNAME (LOCALE_SLOCALIZEDLANGUAGENAME)
value LOCALE_SLANGUAGE (LOCALE_SLOCALIZEDDISPLAYNAME)
value LOCALE_SNATIVECTRYNAME (LOCALE_SNATIVECOUNTRYNAME)
value LOCALE_SNATIVELANGNAME (LOCALE_SNATIVELANGUAGENAME)
value LOCALE_UNASSIGNED_LCID (LOCALE_CUSTOM_UNSPECIFIED)
value LOCK_ELEMENT (0)
value LOGPIXELSX (88)
value LOGPIXELSY (90)
value LONG_MAX (2147483647L)
value LPCPROPSHEETHEADER (LPCPROPSHEETHEADERA)
value LPCPROPSHEETPAGE (LPCPROPSHEETPAGEA)
value LPCPROPSHEETPAGE_LATEST (LPCPROPSHEETPAGEA_LATEST)
value LPD_TYPE_COLORINDEX (1)
value LPD_TYPE_RGBA (0)
value LPFNPSPCALLBACK (LPFNPSPCALLBACKA)
value LPOCNCONNPROC (LPOCNCONNPROCA)
value LPOINET (LPIINTERNET)
value LPOINETBINDINFO (LPIINTERNETBINDINFO)
value LPOINETPRIORITY (LPIINTERNETPRIORITY)
value LPOINETPROTOCOL (LPIINTERNETPROTOCOL)
value LPOINETPROTOCOLEX (LPIINTERNETPROTOCOLEX)
value LPOINETPROTOCOLINFO (LPIINTERNETPROTOCOLINFO)
value LPOINETPROTOCOLROOT (LPIINTERNETPROTOCOLROOT)
value LPOINETPROTOCOLSINK (LPIINTERNETPROTOCOLSINK)
value LPOINETPROTOCOLSINKSTACKABLE (LPIINTERNETPROTOCOLSINKSTACKABLE)
value LPOINETSESSION (LPIINTERNETSESSION)
value LPOINETTHREADSWITCH (LPIINTERNETTHREADSWITCH)
value LPOPENCARDNAMEA_EX (LPOPENCARDNAME_EXA)
value LPOPENCARDNAMEW_EX (LPOPENCARDNAME_EXW)
value LPOPENCARDNAME_A (LPOPENCARDNAMEA)
value LPOPENCARDNAME_W (LPOPENCARDNAMEW)
value LPPROPSHEETHEADER (LPPROPSHEETHEADERA)
value LPPROPSHEETPAGE (LPPROPSHEETPAGEA)
value LPPROPSHEETPAGE_LATEST (LPPROPSHEETPAGEA_LATEST)
value LPSCARD_READERSTATE_A (LPSCARD_READERSTATEA)
value LPSCARD_READERSTATE_W (LPSCARD_READERSTATEW)
value LPSERVICE_MAIN_FUNCTION (LPSERVICE_MAIN_FUNCTIONA)
value LPWSAEVENT (LPHANDLE)
value LSFW_LOCK (1)
value LSFW_UNLOCK (2)
value LTGRAY_BRUSH (1)
value MAC_CHARSET (77)
value MAKEINTRESOURCE (MAKEINTRESOURCEA)
value MARKPARITY (3)
value MARSHALINTERFACE_MIN (500)
value MAXERRORLENGTH (256)
value MAXGETHOSTSTRUCT (1024)
value MAXIMUM_ATTR_STRING_LENGTH (32)
value MAXIMUM_PROCESSORS (MAXIMUM_PROC_PER_GROUP)
value MAXIMUM_PROC_PER_GROUP (64)
value MAXIMUM_SMARTCARD_READERS (10)
value MAXIMUM_SUSPEND_COUNT (MAXCHAR)
value MAXIMUM_WAIT_OBJECTS (64)
value MAXLOGICALLOGNAMESIZE (256)
value MAXPNAMELEN (32)
value MAXPROPPAGES (100)
value MAXSTRETCHBLTMODE (4)
value MAXUIDLEN (64)
value MAX_ACL_REVISION (ACL_REVISION4)
value MAX_COMPUTERNAME_LENGTH (15)
value MAX_DEFAULTCHAR (2)
value MAX_FW_BUCKET_ID_LENGTH (132)
value MAX_HW_COUNTERS (16)
value MAX_INTERFACE_CODES (8)
value MAX_JOYSTICKOEMVXDNAME (260)
value MAX_LANA (254)
value MAX_LEADBYTES (12)
value MAX_LOGICALDPIOVERRIDE (2)
value MAX_MONITORS (4)
value MAX_NUM_REASONS (256)
value MAX_PATH (260)
value MAX_PRIORITY (99)
value MAX_PROFILE_LEN (80)
value MAX_PROTOCOL_CHAIN (7)
value MAX_REASON_BUGID_LEN (32)
value MAX_REASON_COMMENT_LEN (512)
value MAX_REASON_DESC_LEN (256)
value MAX_REASON_NAME_LEN (64)
value MAX_RESOURCEMANAGER_DESCRIPTION_LENGTH (64)
value MAX_SID_SIZE (256)
value MAX_SIZE_SECURITY_ID (512)
value MAX_STR_BLOCKREASON (256)
value MAX_TOUCH_COUNT (256)
value MAX_TOUCH_PREDICTION_FILTER_TAPS (3)
value MAX_TRANSACTION_DESCRIPTION_LENGTH (64)
value MAX_VOLUME_ID_SIZE (36)
value MAX_VOLUME_TEMPLATE_SIZE (40)
value MA_ACTIVATE (1)
value MA_ACTIVATEANDEAT (2)
value MA_NOACTIVATE (3)
value MA_NOACTIVATEANDEAT (4)
value MB_ICONERROR (MB_ICONHAND)
value MB_ICONINFORMATION (MB_ICONASTERISK)
value MB_ICONSTOP (MB_ICONHAND)
value MB_ICONWARNING (MB_ICONEXCLAMATION)
value MB_LEN_MAX (5)
value MCIERR_BASE (256)
value MCI_CD_OFFSET (1088)
value MCI_DEVTYPE_ANIMATION (519)
value MCI_DEVTYPE_CD_AUDIO (516)
value MCI_DEVTYPE_DAT (517)
value MCI_DEVTYPE_DIGITAL_VIDEO (520)
value MCI_DEVTYPE_FIRST (MCI_DEVTYPE_VCR)
value MCI_DEVTYPE_LAST (MCI_DEVTYPE_SEQUENCER)
value MCI_DEVTYPE_OTHER (521)
value MCI_DEVTYPE_OVERLAY (515)
value MCI_DEVTYPE_SCANNER (518)
value MCI_DEVTYPE_SEQUENCER (523)
value MCI_DEVTYPE_VCR (513)
value MCI_DEVTYPE_VIDEODISC (514)
value MCI_DEVTYPE_WAVEFORM_AUDIO (522)
value MCI_FIRST (DRV_MCI_FIRST)
value MCI_FORMAT_BYTES (8)
value MCI_FORMAT_FRAMES (3)
value MCI_FORMAT_HMS (1)
value MCI_FORMAT_MILLISECONDS (0)
value MCI_FORMAT_MSF (2)
value MCI_FORMAT_SAMPLES (9)
value MCI_FORMAT_TMSF (10)
value MCI_SEQ_MAPPER (65535)
value MCI_SEQ_NONE (65533)
value MCI_SEQ_OFFSET (1216)
value MCI_STRING_OFFSET (512)
value MCI_VD_OFFSET (1024)
value MCI_WAVE_OFFSET (1152)
value MDM_PIAFS_INCOMING (0)
value MDM_PIAFS_OUTGOING (1)
value MDM_SHIFT_BEARERMODE (12)
value MDM_SHIFT_EXTENDEDINFO (MDM_SHIFT_BEARERMODE)
value MDM_SHIFT_PROTOCOLDATA (20)
value MDM_SHIFT_PROTOCOLID (16)
value MDM_SHIFT_PROTOCOLINFO (MDM_SHIFT_PROTOCOLID)
value MEMBERID_NIL (DISPID_UNKNOWN)
value MEMORY_ALLOCATION_ALIGNMENT (16)
value MEMORY_PRIORITY_BELOW_NORMAL (4)
value MEMORY_PRIORITY_LOW (2)
value MEMORY_PRIORITY_LOWEST (0)
value MEMORY_PRIORITY_MEDIUM (3)
value MEMORY_PRIORITY_NORMAL (5)
value MEMORY_PRIORITY_VERY_LOW (1)
value MEM_EXTENDED_PARAMETER_NUMA_NODE_MANDATORY (MINLONG64)
value MEM_EXTENDED_PARAMETER_TYPE_BITS (8)
value METAFILE_DRIVER (2049)
value METHOD_BUFFERED (0)
value METHOD_DIRECT_FROM_HARDWARE (METHOD_OUT_DIRECT)
value METHOD_DIRECT_TO_HARDWARE (METHOD_IN_DIRECT)
value METHOD_IN_DIRECT (1)
value METHOD_NEITHER (3)
value METHOD_OUT_DIRECT (2)
value MFCOMMENT (15)
value MFS_CHECKED (MF_CHECKED)
value MFS_DEFAULT (MF_DEFAULT)
value MFS_DISABLED (MFS_GRAYED)
value MFS_ENABLED (MF_ENABLED)
value MFS_HILITE (MF_HILITE)
value MFS_UNCHECKED (MF_UNCHECKED)
value MFS_UNHILITE (MF_UNHILITE)
value MFT_BITMAP (MF_BITMAP)
value MFT_MENUBARBREAK (MF_MENUBARBREAK)
value MFT_MENUBREAK (MF_MENUBREAK)
value MFT_OWNERDRAW (MF_OWNERDRAW)
value MFT_RIGHTJUSTIFY (MF_RIGHTJUSTIFY)
value MFT_SEPARATOR (MF_SEPARATOR)
value MFT_STRING (MF_STRING)
value MH_CLEANUP (4)
value MH_CREATE (1)
value MH_DELETE (3)
value MH_KEEP (2)
value MICROSOFT_WINBASE_H_DEFINE_INTERLOCKED_CPLUSPLUS_OVERLOADS (0)
value MICROSOFT_WINDOWS_WINBASE_H_DEFINE_INTERLOCKED_CPLUSPLUS_OVERLOADS (1)
value MIDIERR_BASE (64)
value MIDIPATCHSIZE (128)
value MIDI_CACHE_ALL (1)
value MIDI_CACHE_BESTFIT (2)
value MIDI_CACHE_QUERY (3)
value MIDI_UNCACHE (4)
value MIM_CLOSE (MM_MIM_CLOSE)
value MIM_DATA (MM_MIM_DATA)
value MIM_ERROR (MM_MIM_ERROR)
value MIM_LONGDATA (MM_MIM_LONGDATA)
value MIM_LONGERROR (MM_MIM_LONGERROR)
value MIM_MOREDATA (MM_MIM_MOREDATA)
value MIM_OPEN (MM_MIM_OPEN)
value MIN_ACL_REVISION (ACL_REVISION2)
value MIN_PRIORITY (1)
value MIXERLINE_TARGETTYPE_AUX (5)
value MIXERLINE_TARGETTYPE_MIDIIN (4)
value MIXERLINE_TARGETTYPE_MIDIOUT (3)
value MIXERLINE_TARGETTYPE_UNDEFINED (0)
value MIXERLINE_TARGETTYPE_WAVEIN (2)
value MIXERLINE_TARGETTYPE_WAVEOUT (1)
value MIXERR_BASE (1024)
value MIXER_LONG_NAME_CHARS (64)
value MIXER_SHORT_NAME_CHARS (16)
value MKSYS_URLMONIKER (6)
value MMIOERR_BASE (256)
value MMIOM_CLOSE (4)
value MMIOM_OPEN (3)
value MMIOM_READ (MMIO_READ)
value MMIOM_RENAME (6)
value MMIOM_SEEK (2)
value MMIOM_WRITE (MMIO_WRITE)
value MMIOM_WRITEFLUSH (5)
value MMIO_DEFAULTBUFFER (8192)
value MMSYSERR_BASE (0)
value MMSYSERR_NOERROR (0)
value MM_ANISOTROPIC (8)
value MM_HIENGLISH (5)
value MM_HIMETRIC (3)
value MM_ISOTROPIC (7)
value MM_LOENGLISH (4)
value MM_LOMETRIC (2)
value MM_MAX (MM_ANISOTROPIC)
value MM_MAX_AXES_NAMELEN (16)
value MM_MAX_FIXEDSCALE (MM_TWIPS)
value MM_MAX_NUMAXES (16)
value MM_MIN (MM_TEXT)
value MM_TEXT (1)
value MM_TWIPS (6)
value MNC_CLOSE (1)
value MNC_EXECUTE (2)
value MNC_IGNORE (0)
value MNC_SELECT (3)
value MND_CONTINUE (0)
value MND_ENDMENU (1)
value MOD_FMSYNTH (4)
value MOD_MAPPER (5)
value MOD_MIDIPORT (1)
value MOD_SQSYNTH (3)
value MOD_SWSYNTH (7)
value MOD_SYNTH (2)
value MOD_WAVETABLE (6)
value MOM_CLOSE (MM_MOM_CLOSE)
value MOM_DONE (MM_MOM_DONE)
value MOM_OPEN (MM_MOM_OPEN)
value MOM_POSITIONCB (MM_MOM_POSITIONCB)
value MONO_FONT (8)
value MOUSETRAILS (39)
value MOUSEWHEEL_ROUTING_FOCUS (0)
value MOUSEWHEEL_ROUTING_HYBRID (1)
value MOUSEWHEEL_ROUTING_MOUSE_POS (2)
value MOUSE_MOVE_ABSOLUTE (1)
value MOUSE_MOVE_RELATIVE (0)
value MSGFLT_ADD (1)
value MSGFLT_REMOVE (2)
value MSGF_DIALOGBOX (0)
value MSGF_MAX (8)
value MSGF_MENU (2)
value MSGF_MESSAGEBOX (1)
value MSGF_NEXTWINDOW (6)
value MSGF_SCROLLBAR (5)
value MSGF_USER (4096)
value MSG_MAXIOVLEN (16)
value MS_DEF_DH_SCHANNEL_PROV (MS_DEF_DH_SCHANNEL_PROV_A)
value MS_DEF_DSS_DH_PROV (MS_DEF_DSS_DH_PROV_A)
value MS_DEF_DSS_PROV (MS_DEF_DSS_PROV_A)
value MS_DEF_PROV (MS_DEF_PROV_A)
value MS_DEF_RSA_SCHANNEL_PROV (MS_DEF_RSA_SCHANNEL_PROV_A)
value MS_DEF_RSA_SIG_PROV (MS_DEF_RSA_SIG_PROV_A)
value MS_ENHANCED_PROV (MS_ENHANCED_PROV_A)
value MS_ENH_DSS_DH_PROV (MS_ENH_DSS_DH_PROV_A)
value MS_ENH_RSA_AES_PROV (MS_ENH_RSA_AES_PROV_A)
value MS_ENH_RSA_AES_PROV_XP (MS_ENH_RSA_AES_PROV_XP_A)
value MS_SCARD_PROV (MS_SCARD_PROV_A)
value MS_STRONG_PROV (MS_STRONG_PROV_A)
value MUI_CALLBACK_ALL_FLAGS (MUI_CALLBACK_FLAG_UPGRADED_INSTALLATION)
value MULTIFILEOPENORD (1537)
value MUTEX_ALL_ACCESS (MUTANT_ALL_ACCESS)
value MUTEX_MODIFY_STATE (MUTANT_QUERY_STATE)
value MWT_IDENTITY (1)
value MWT_LEFTMULTIPLY (2)
value MWT_MAX (MWT_RIGHTMULTIPLY)
value MWT_MIN (MWT_IDENTITY)
value MWT_RIGHTMULTIPLY (3)
value NCBNAMSZ (16)
value NCRYPTBUFFER_ATTESTATIONSTATEMENT_BLOB (51)
value NCRYPTBUFFER_ATTESTATION_CLAIM_CHALLENGE_REQUIRED (53)
value NCRYPTBUFFER_ATTESTATION_CLAIM_TYPE (52)
value NCRYPTBUFFER_CERT_BLOB (47)
value NCRYPTBUFFER_CLAIM_IDBINDING_NONCE (48)
value NCRYPTBUFFER_CLAIM_KEYATTESTATION_NONCE (49)
value NCRYPTBUFFER_DATA (1)
value NCRYPTBUFFER_ECC_CURVE_NAME (60)
value NCRYPTBUFFER_ECC_PARAMETERS (61)
value NCRYPTBUFFER_EMPTY (0)
value NCRYPTBUFFER_KEY_PROPERTY_FLAGS (50)
value NCRYPTBUFFER_PKCS_ALG_ID (43)
value NCRYPTBUFFER_PKCS_ALG_OID (41)
value NCRYPTBUFFER_PKCS_ALG_PARAM (42)
value NCRYPTBUFFER_PKCS_ATTRS (44)
value NCRYPTBUFFER_PKCS_KEY_NAME (45)
value NCRYPTBUFFER_PKCS_OID (40)
value NCRYPTBUFFER_PKCS_SECRET (46)
value NCRYPTBUFFER_PROTECTION_DESCRIPTOR_STRING (3)
value NCRYPTBUFFER_PROTECTION_FLAGS (4)
value NCRYPTBUFFER_SSL_CLEAR_KEY (23)
value NCRYPTBUFFER_SSL_CLIENT_RANDOM (20)
value NCRYPTBUFFER_SSL_HIGHEST_VERSION (22)
value NCRYPTBUFFER_SSL_KEY_ARG_DATA (24)
value NCRYPTBUFFER_SSL_SERVER_RANDOM (21)
value NCRYPTBUFFER_SSL_SESSION_HASH (25)
value NCRYPTBUFFER_TPM_PLATFORM_CLAIM_NONCE (81)
value NCRYPTBUFFER_TPM_PLATFORM_CLAIM_PCR_MASK (80)
value NCRYPTBUFFER_TPM_PLATFORM_CLAIM_STATIC_CREATE (82)
value NCRYPTBUFFER_TPM_SEAL_NO_DA_PROTECTION (73)
value NCRYPTBUFFER_TPM_SEAL_PASSWORD (70)
value NCRYPTBUFFER_TPM_SEAL_POLICYINFO (71)
value NCRYPTBUFFER_TPM_SEAL_TICKET (72)
value NCRYPTBUFFER_VERSION (0)
value NCRYPTBUFFER_VSM_KEY_ATTESTATION_CLAIM_RESTRICTIONS (54)
value NCRYPT_AES_ALGORITHM (BCRYPT_AES_ALGORITHM)
value NCRYPT_AES_ALGORITHM_GROUP (NCRYPT_AES_ALGORITHM)
value NCRYPT_ALTERNATE_KEY_STORAGE_LOCATION_PROPERTY (NCRYPT_PCP_ALTERNATE_KEY_STORAGE_LOCATION_PROPERTY)
value NCRYPT_ASYMMETRIC_ENCRYPTION_INTERFACE (BCRYPT_ASYMMETRIC_ENCRYPTION_INTERFACE)
value NCRYPT_ASYMMETRIC_ENCRYPTION_OPERATION (BCRYPT_ASYMMETRIC_ENCRYPTION_OPERATION)
value NCRYPT_CAPI_KDF_ALGORITHM (BCRYPT_CAPI_KDF_ALGORITHM)
value NCRYPT_CHANGEPASSWORD_PROPERTY (NCRYPT_PCP_CHANGEPASSWORD_PROPERTY)
value NCRYPT_CIPHER_INTERFACE (BCRYPT_CIPHER_INTERFACE)
value NCRYPT_CIPHER_OPERATION (BCRYPT_CIPHER_OPERATION)
value NCRYPT_DESX_ALGORITHM (BCRYPT_DESX_ALGORITHM)
value NCRYPT_DES_ALGORITHM (BCRYPT_DES_ALGORITHM)
value NCRYPT_DH_ALGORITHM (BCRYPT_DH_ALGORITHM)
value NCRYPT_DH_ALGORITHM_GROUP (NCRYPT_DH_ALGORITHM)
value NCRYPT_DH_PARAMETERS_PROPERTY (BCRYPT_DH_PARAMETERS)
value NCRYPT_DSA_ALGORITHM (BCRYPT_DSA_ALGORITHM)
value NCRYPT_DSA_ALGORITHM_GROUP (NCRYPT_DSA_ALGORITHM)
value NCRYPT_ECC_CURVE_NAME_LIST_PROPERTY (BCRYPT_ECC_CURVE_NAME_LIST)
value NCRYPT_ECC_CURVE_NAME_PROPERTY (BCRYPT_ECC_CURVE_NAME)
value NCRYPT_ECC_PARAMETERS_PROPERTY (BCRYPT_ECC_PARAMETERS)
value NCRYPT_ECDH_ALGORITHM (BCRYPT_ECDH_ALGORITHM)
value NCRYPT_ECDSA_ALGORITHM (BCRYPT_ECDSA_ALGORITHM)
value NCRYPT_EXPORTED_ISOLATED_KEY_HEADER_CURRENT_VERSION (NCRYPT_EXPORTED_ISOLATED_KEY_HEADER_V0)
value NCRYPT_HASH_INTERFACE (BCRYPT_HASH_INTERFACE)
value NCRYPT_HASH_OPERATION (BCRYPT_HASH_OPERATION)
value NCRYPT_INITIALIZATION_VECTOR (BCRYPT_INITIALIZATION_VECTOR)
value NCRYPT_ISOLATED_KEY_ATTESTED_ATTRIBUTES_CURRENT_VERSION (NCRYPT_ISOLATED_KEY_ATTESTED_ATTRIBUTES_V0)
value NCRYPT_KEY_ACCESS_POLICY_VERSION (1)
value NCRYPT_KEY_DERIVATION_INTERFACE (BCRYPT_KEY_DERIVATION_INTERFACE)
value NCRYPT_KEY_DERIVATION_OPERATION (BCRYPT_KEY_DERIVATION_OPERATION)
value NCRYPT_MAX_ALG_ID_LENGTH (512)
value NCRYPT_MAX_KEY_NAME_LENGTH (512)
value NCRYPT_MAX_PROPERTY_NAME (64)
value NCRYPT_NO_KEY_VALIDATION (BCRYPT_NO_KEY_VALIDATION)
value NCRYPT_PIN_CACHE_APPLICATION_TICKET_BYTE_LENGTH (90)
value NCRYPT_PIN_CACHE_PIN_BYTE_LENGTH (90)
value NCRYPT_PUBLIC_LENGTH_PROPERTY (BCRYPT_PUBLIC_KEY_LENGTH)
value NCRYPT_RNG_OPERATION (BCRYPT_RNG_OPERATION)
value NCRYPT_RSA_ALGORITHM (BCRYPT_RSA_ALGORITHM)
value NCRYPT_RSA_ALGORITHM_GROUP (NCRYPT_RSA_ALGORITHM)
value NCRYPT_RSA_SIGN_ALGORITHM (BCRYPT_RSA_SIGN_ALGORITHM)
value NCRYPT_SECRET_AGREEMENT_INTERFACE (BCRYPT_SECRET_AGREEMENT_INTERFACE)
value NCRYPT_SECRET_AGREEMENT_OPERATION (BCRYPT_SECRET_AGREEMENT_OPERATION)
value NCRYPT_SIGNATURE_INTERFACE (BCRYPT_SIGNATURE_INTERFACE)
value NCRYPT_SIGNATURE_LENGTH_PROPERTY (BCRYPT_SIGNATURE_LENGTH)
value NCRYPT_SIGNATURE_OPERATION (BCRYPT_SIGNATURE_OPERATION)
value NCRYPT_TPM_PLATFORM_ATTESTATION_STATEMENT_CURRENT_VERSION (NCRYPT_TPM_PLATFORM_ATTESTATION_STATEMENT_V0)
value NCRYPT_VSM_KEY_ATTESTATION_CLAIM_RESTRICTIONS_CURRENT_VERSION (NCRYPT_VSM_KEY_ATTESTATION_CLAIM_RESTRICTIONS_V0)
value NCRYPT_VSM_KEY_ATTESTATION_STATEMENT_CURRENT_VERSION (NCRYPT_VSM_KEY_ATTESTATION_STATEMENT_V0)
value NDR_LOCAL_ENDIAN (NDR_LITTLE_ENDIAN)
value NETPROPERTY_PERSISTENT (1)
value NEWFILEOPENORD (1547)
value NEWFORMATDLGWITHLINK (1591)
value NEWFRAME (1)
value NEWTRANSPARENT (3)
value NEXTBAND (3)
value NFR_ANSI (1)
value NFR_UNICODE (2)
value NF_QUERY (3)
value NF_REQUERY (4)
value NI_MAXHOST (1025)
value NI_MAXSERV (32)
value NOERROR (0)
value NONANTIALIASED_QUALITY (3)
value NOPARITY (0)
value NOTIFYICON_VERSION (3)
value NO_ADDRESS (WSANO_ADDRESS)
value NO_DATA (WSANO_DATA)
value NO_ERROR (0cL)
value NO_PRIORITY (0)
value NO_RECOVERY (WSANO_RECOVERY)
value NTAPI_INLINE (NTAPI)
value NTDDI_LONGHORN (NTDDI_VISTA)
value NTDDI_VERSION (WDK_NTDDI_VERSION)
value NTDDI_VISTA (NTDDI_WIN6)
value NTE_OP_OK (0)
value NTSYSAPI (DECLSPEC_IMPORT)
value NTSYSCALLAPI (DECLSPEC_IMPORT)
value NULLREGION (1)
value NULL_BRUSH (5)
value NULL_PEN (8)
value NUMBRUSHES (16)
value NUMCOLORS (24)
value NUMFONTS (22)
value NUMMARKERS (20)
value NUMPENS (18)
value NUMRESERVED (106)
value NUM_DISCHARGE_POLICIES (4)
value N_BTSHFT (4)
value N_TSHIFT (2)
value OBJ_BITMAP (7)
value OBJ_BRUSH (2)
value OBJ_COLORSPACE (14)
value OBJ_DC (3)
value OBJ_ENHMETADC (12)
value OBJ_ENHMETAFILE (13)
value OBJ_EXTPEN (11)
value OBJ_FONT (6)
value OBJ_MEMDC (10)
value OBJ_METADC (4)
value OBJ_METAFILE (9)
value OBJ_PAL (5)
value OBJ_PEN (1)
value OBJ_REGION (8)
value OCSP_BASIC_BY_KEY_RESPONDER_ID (2)
value OCSP_BASIC_BY_NAME_RESPONDER_ID (1)
value OCSP_BASIC_GOOD_CERT_STATUS (0)
value OCSP_BASIC_REVOKED_CERT_STATUS (1)
value OCSP_BASIC_UNKNOWN_CERT_STATUS (2)
value OCSP_INTERNAL_ERROR_RESPONSE (2)
value OCSP_MALFORMED_REQUEST_RESPONSE (1)
value OCSP_SIG_REQUIRED_RESPONSE (5)
value OCSP_SUCCESSFUL_RESPONSE (0)
value OCSP_TRY_LATER_RESPONSE (3)
value OCSP_UNAUTHORIZED_RESPONSE (6)
value ODDPARITY (1)
value ODT_BUTTON (4)
value ODT_COMBOBOX (3)
value ODT_LISTBOX (2)
value ODT_MENU (1)
value ODT_STATIC (5)
value OEM_CHARSET (255)
value OEM_FIXED_FONT (10)
value OFN_SHAREFALLTHROUGH (2)
value OFN_SHARENOWARN (1)
value OFN_SHAREWARN (0)
value OFS_MAXPATHNAME (128)
value OLDFONTENUMPROC (OLDFONTENUMPROCA)
value ONESTOPBIT (0)
value OPAQUE (2)
value OPENCARDNAMEA_EX (OPENCARDNAME_EXA)
value OPENCARDNAMEW_EX (OPENCARDNAME_EXW)
value OPENCARDNAME_A (OPENCARDNAMEA)
value OPENCARDNAME_W (OPENCARDNAMEW)
value OPENCHANNEL (4110)
value OPEN_ALWAYS (4)
value OPEN_EXISTING (3)
value OPERATION_API_VERSION (1)
value ORD_LANGDRIVER (1)
value OR_INVALID_OID (1911L)
value OR_INVALID_OXID (1910L)
value OR_INVALID_SET (1912L)
value OUTPUT_DEBUG_STRING_EVENT (8)
value OUT_CHARACTER_PRECIS (2)
value OUT_DEFAULT_PRECIS (0)
value OUT_DEVICE_PRECIS (5)
value OUT_OUTLINE_PRECIS (8)
value OUT_PS_ONLY_PRECIS (10)
value OUT_RASTER_PRECIS (6)
value OUT_SCREEN_OUTLINE_PRECIS (9)
value OUT_STRING_PRECIS (1)
value OUT_STROKE_PRECIS (3)
value OUT_TT_ONLY_PRECIS (7)
value OUT_TT_PRECIS (4)
value O_APPEND (_O_APPEND)
value O_BINARY (_O_BINARY)
value O_CREAT (_O_CREAT)
value O_EXCL (_O_EXCL)
value O_NOINHERIT (_O_NOINHERIT)
value O_RANDOM (_O_RANDOM)
value O_RAW (_O_BINARY)
value O_RDONLY (_O_RDONLY)
value O_RDWR (_O_RDWR)
value O_SEQUENTIAL (_O_SEQUENTIAL)
value O_TEMPORARY (_O_TEMPORARY)
value O_TEXT (_O_TEXT)
value O_TRUNC (_O_TRUNC)
value O_WRONLY (_O_WRONLY)
value PAGESETUPDLGORD (1546)
value PAGESETUPDLGORDMOTIF (1550)
value PANOSE_COUNT (10)
value PAN_ANY (0)
value PAN_ARMSTYLE_INDEX (6)
value PAN_BENT_ARMS_DOUBLE_SERIF (11)
value PAN_BENT_ARMS_HORZ (7)
value PAN_BENT_ARMS_SINGLE_SERIF (10)
value PAN_BENT_ARMS_VERT (9)
value PAN_BENT_ARMS_WEDGE (8)
value PAN_CONTRAST_HIGH (8)
value PAN_CONTRAST_INDEX (4)
value PAN_CONTRAST_LOW (4)
value PAN_CONTRAST_MEDIUM (6)
value PAN_CONTRAST_MEDIUM_HIGH (7)
value PAN_CONTRAST_MEDIUM_LOW (5)
value PAN_CONTRAST_NONE (2)
value PAN_CONTRAST_VERY_HIGH (9)
value PAN_CONTRAST_VERY_LOW (3)
value PAN_CULTURE_LATIN (0)
value PAN_FAMILYTYPE_INDEX (0)
value PAN_FAMILY_DECORATIVE (4)
value PAN_FAMILY_PICTORIAL (5)
value PAN_FAMILY_SCRIPT (3)
value PAN_FAMILY_TEXT_DISPLAY (2)
value PAN_LETTERFORM_INDEX (7)
value PAN_LETT_NORMAL_BOXED (4)
value PAN_LETT_NORMAL_CONTACT (2)
value PAN_LETT_NORMAL_FLATTENED (5)
value PAN_LETT_NORMAL_OFF_CENTER (7)
value PAN_LETT_NORMAL_ROUNDED (6)
value PAN_LETT_NORMAL_SQUARE (8)
value PAN_LETT_NORMAL_WEIGHTED (3)
value PAN_LETT_OBLIQUE_BOXED (11)
value PAN_LETT_OBLIQUE_CONTACT (9)
value PAN_LETT_OBLIQUE_FLATTENED (12)
value PAN_LETT_OBLIQUE_OFF_CENTER (14)
value PAN_LETT_OBLIQUE_ROUNDED (13)
value PAN_LETT_OBLIQUE_SQUARE (15)
value PAN_LETT_OBLIQUE_WEIGHTED (10)
value PAN_MIDLINE_CONSTANT_POINTED (9)
value PAN_MIDLINE_CONSTANT_SERIFED (10)
value PAN_MIDLINE_CONSTANT_TRIMMED (8)
value PAN_MIDLINE_HIGH_POINTED (6)
value PAN_MIDLINE_HIGH_SERIFED (7)
value PAN_MIDLINE_HIGH_TRIMMED (5)
value PAN_MIDLINE_INDEX (8)
value PAN_MIDLINE_LOW_POINTED (12)
value PAN_MIDLINE_LOW_SERIFED (13)
value PAN_MIDLINE_LOW_TRIMMED (11)
value PAN_MIDLINE_STANDARD_POINTED (3)
value PAN_MIDLINE_STANDARD_SERIFED (4)
value PAN_MIDLINE_STANDARD_TRIMMED (2)
value PAN_NO_FIT (1)
value PAN_PROPORTION_INDEX (3)
value PAN_PROP_CONDENSED (6)
value PAN_PROP_EVEN_WIDTH (4)
value PAN_PROP_EXPANDED (5)
value PAN_PROP_MODERN (3)
value PAN_PROP_MONOSPACED (9)
value PAN_PROP_OLD_STYLE (2)
value PAN_PROP_VERY_CONDENSED (8)
value PAN_PROP_VERY_EXPANDED (7)
value PAN_SERIFSTYLE_INDEX (1)
value PAN_SERIF_BONE (8)
value PAN_SERIF_COVE (2)
value PAN_SERIF_EXAGGERATED (9)
value PAN_SERIF_FLARED (14)
value PAN_SERIF_NORMAL_SANS (11)
value PAN_SERIF_OBTUSE_COVE (3)
value PAN_SERIF_OBTUSE_SANS (12)
value PAN_SERIF_OBTUSE_SQUARE_COVE (5)
value PAN_SERIF_PERP_SANS (13)
value PAN_SERIF_ROUNDED (15)
value PAN_SERIF_SQUARE (6)
value PAN_SERIF_SQUARE_COVE (4)
value PAN_SERIF_THIN (7)
value PAN_SERIF_TRIANGLE (10)
value PAN_STRAIGHT_ARMS_DOUBLE_SERIF (6)
value PAN_STRAIGHT_ARMS_HORZ (2)
value PAN_STRAIGHT_ARMS_SINGLE_SERIF (5)
value PAN_STRAIGHT_ARMS_VERT (4)
value PAN_STRAIGHT_ARMS_WEDGE (3)
value PAN_STROKEVARIATION_INDEX (5)
value PAN_STROKE_GRADUAL_DIAG (2)
value PAN_STROKE_GRADUAL_HORZ (5)
value PAN_STROKE_GRADUAL_TRAN (3)
value PAN_STROKE_GRADUAL_VERT (4)
value PAN_STROKE_INSTANT_VERT (8)
value PAN_STROKE_RAPID_HORZ (7)
value PAN_STROKE_RAPID_VERT (6)
value PAN_WEIGHT_BLACK (10)
value PAN_WEIGHT_BOLD (8)
value PAN_WEIGHT_BOOK (5)
value PAN_WEIGHT_DEMI (7)
value PAN_WEIGHT_HEAVY (9)
value PAN_WEIGHT_INDEX (2)
value PAN_WEIGHT_LIGHT (3)
value PAN_WEIGHT_MEDIUM (6)
value PAN_WEIGHT_NORD (11)
value PAN_WEIGHT_THIN (4)
value PAN_WEIGHT_VERY_LIGHT (2)
value PAN_XHEIGHT_CONSTANT_LARGE (4)
value PAN_XHEIGHT_CONSTANT_SMALL (2)
value PAN_XHEIGHT_CONSTANT_STD (3)
value PAN_XHEIGHT_DUCKING_LARGE (7)
value PAN_XHEIGHT_DUCKING_SMALL (5)
value PAN_XHEIGHT_DUCKING_STD (6)
value PAN_XHEIGHT_INDEX (9)
value PARKING_TOPOLOGY_POLICY_DISABLED (0)
value PARKING_TOPOLOGY_POLICY_ROUNDROBIN (1)
value PARKING_TOPOLOGY_POLICY_SEQUENTIAL (2)
value PARSE_DECODE (PARSE_DECODE_IS_ESCAPE)
value PARSE_ENCODE (PARSE_ENCODE_IS_UNESCAPE)
value PASSEMBLY_DLL_REDIRECTION_DETAILED_INFORMATION (PASSEMBLY_FILE_DETAILED_INFORMATION)
value PASSIVE_LEVEL (0)
value PASSTHROUGH (19)
value PA_ACTIVATE (MA_ACTIVATE)
value PA_NOACTIVATE (MA_NOACTIVATE)
value PCASSEMBLY_DLL_REDIRECTION_DETAILED_INFORMATION (PCASSEMBLY_FILE_DETAILED_INFORMATION)
value PC_INTERIORS (128)
value PC_NONE (0)
value PC_PATHS (512)
value PC_POLYGON (1)
value PC_POLYPOLYGON (256)
value PC_RECTANGLE (2)
value PC_SCANLINE (8)
value PC_STYLED (32)
value PC_TRAPEZOID (4)
value PC_WIDE (16)
value PC_WIDESTYLED (64)
value PC_WINDPOLYGON (4)
value PDEVICESIZE (26)
value PD_RESULT_APPLY (2)
value PD_RESULT_CANCEL (0)
value PD_RESULT_PRINT (1)
value PEERDIST_ERROR_ALREADY_COMPLETED (4060L)
value PEERDIST_ERROR_ALREADY_EXISTS (4058L)
value PEERDIST_ERROR_ALREADY_INITIALIZED (4055L)
value PEERDIST_ERROR_CANNOT_PARSE_CONTENTINFO (4051L)
value PEERDIST_ERROR_CONTENTINFO_VERSION_UNSUPPORTED (4050L)
value PEERDIST_ERROR_INVALIDATED (4057L)
value PEERDIST_ERROR_INVALID_CONFIGURATION (4063L)
value PEERDIST_ERROR_MISSING_DATA (4052L)
value PEERDIST_ERROR_NOT_INITIALIZED (4054L)
value PEERDIST_ERROR_NOT_LICENSED (4064L)
value PEERDIST_ERROR_NO_MORE (4053L)
value PEERDIST_ERROR_OPERATION_NOTFOUND (4059L)
value PEERDIST_ERROR_OUT_OF_BOUNDS (4061L)
value PEERDIST_ERROR_SERVICE_UNAVAILABLE (4065L)
value PEERDIST_ERROR_SHUTDOWN_IN_PROGRESS (4056L)
value PEERDIST_ERROR_TRUST_FAILURE (4066L)
value PEERDIST_ERROR_VERSION_UNSUPPORTED (4062L)
value PERFORMANCE_DATA_VERSION (1)
value PERFSTATE_POLICY_CHANGE_DECREASE_MAX (PERFSTATE_POLICY_CHANGE_ROCKET)
value PERFSTATE_POLICY_CHANGE_IDEAL (0)
value PERFSTATE_POLICY_CHANGE_IDEAL_AGGRESSIVE (3)
value PERFSTATE_POLICY_CHANGE_INCREASE_MAX (PERFSTATE_POLICY_CHANGE_IDEAL_AGGRESSIVE)
value PERFSTATE_POLICY_CHANGE_ROCKET (2)
value PERFSTATE_POLICY_CHANGE_SINGLE (1)
value PERF_DATA_REVISION (1)
value PERF_DATA_VERSION (1)
value PERF_DETAIL_ADVANCED (200)
value PERF_DETAIL_EXPERT (300)
value PERF_DETAIL_NOVICE (100)
value PERF_DETAIL_WIZARD (400)
value PERF_PRECISION_TIMESTAMP (PERF_LARGE_RAW_BASE)
value PFD_MAIN_PLANE (0)
value PFD_OVERLAY_PLANE (1)
value PFD_TYPE_COLORINDEX (1)
value PFD_TYPE_RGBA (0)
value PFORCEINLINE (FORCEINLINE)
value PF_ALPHA_BYTE_INSTRUCTIONS (5)
value PF_APPLETALK (AF_APPLETALK)
value PF_ARM_DIVIDE_INSTRUCTION_AVAILABLE (24)
value PF_ARM_EXTERNAL_CACHE_AVAILABLE (26)
value PF_ARM_FMAC_INSTRUCTIONS_AVAILABLE (27)
value PF_ARM_NEON_INSTRUCTIONS_AVAILABLE (19)
value PF_ATM (AF_ATM)
value PF_AVX_INSTRUCTIONS_AVAILABLE (39)
value PF_BAN (AF_BAN)
value PF_BTH (AF_BTH)
value PF_CCITT (AF_CCITT)
value PF_CHANNELS_ENABLED (16)
value PF_CHAOS (AF_CHAOS)
value PF_COMPARE_EXCHANGE_DOUBLE (2)
value PF_DATAKIT (AF_DATAKIT)
value PF_DLI (AF_DLI)
value PF_ECMA (AF_ECMA)
value PF_ERMS_AVAILABLE (42)
value PF_FASTFAIL_AVAILABLE (23)
value PF_FIREFOX (AF_FIREFOX)
value PF_FLOATING_POINT_EMULATED (1)
value PF_FLOATING_POINT_PRECISION_ERRATA (0)
value PF_HYLINK (AF_HYLINK)
value PF_IMPLINK (AF_IMPLINK)
value PF_INET (AF_INET)
value PF_IPX (AF_IPX)
value PF_ISO (AF_ISO)
value PF_LAT (AF_LAT)
value PF_MAX (AF_MAX)
value PF_MMX_INSTRUCTIONS_AVAILABLE (3)
value PF_MONITORX_INSTRUCTION_AVAILABLE (35)
value PF_NON_TEMPORAL_LEVEL_ALL (_MM_HINT_NTA)
value PF_NS (AF_NS)
value PF_NX_ENABLED (12)
value PF_OSI (AF_OSI)
value PF_PAE_ENABLED (9)
value PF_PUP (AF_PUP)
value PF_RDPID_INSTRUCTION_AVAILABLE (33)
value PF_RDRAND_INSTRUCTION_AVAILABLE (28)
value PF_RDTSCP_INSTRUCTION_AVAILABLE (32)
value PF_RDTSC_INSTRUCTION_AVAILABLE (8)
value PF_RDWRFSGSBASE_AVAILABLE (22)
value PF_SECOND_LEVEL_ADDRESS_TRANSLATION (20)
value PF_SNA (AF_SNA)
value PF_SSE_DAZ_MODE_AVAILABLE (11)
value PF_UNIX (AF_UNIX)
value PF_UNSPEC (AF_UNSPEC)
value PF_VIRT_FIRMWARE_ENABLED (21)
value PF_VOICEVIEW (AF_VOICEVIEW)
value PF_XMMI_INSTRUCTIONS_AVAILABLE (6)
value PF_XSAVE_ENABLED (17)
value PGET_MODULE_HANDLE_EX (PGET_MODULE_HANDLE_EXA)
value PHYSICALHEIGHT (111)
value PHYSICALOFFSETX (112)
value PHYSICALOFFSETY (113)
value PHYSICALWIDTH (110)
value PIPE_UNLIMITED_INSTANCES (255)
value PI_DOCFILECLSIDLOOKUP (PI_CLSIDLOOKUP)
value PKCS_RSA_SSA_PSS_TRAILER_FIELD_BC (1)
value PLANES (14)
value PME_CURRENT_VERSION (1)
value POINTER_DEVICE_PRODUCT_STRING_MAX (520)
value POLICY_SHOWREASONUI_ALWAYS (1)
value POLICY_SHOWREASONUI_NEVER (0)
value POLICY_SHOWREASONUI_SERVERONLY (3)
value POLICY_SHOWREASONUI_WORKSTATIONONLY (2)
value POLYFILL_LAST (2)
value POLYGONALCAPS (32)
value POPENCARDNAMEA_EX (POPENCARDNAME_EXA)
value POPENCARDNAMEW_EX (POPENCARDNAME_EXW)
value POPENCARDNAME_A (POPENCARDNAMEA)
value POPENCARDNAME_W (POPENCARDNAMEW)
value PORT_STATUS_DOOR_OPEN (7)
value PORT_STATUS_NO_TONER (6)
value PORT_STATUS_OFFLINE (1)
value PORT_STATUS_OUTPUT_BIN_FULL (4)
value PORT_STATUS_OUT_OF_MEMORY (9)
value PORT_STATUS_PAPER_JAM (2)
value PORT_STATUS_PAPER_OUT (3)
value PORT_STATUS_PAPER_PROBLEM (5)
value PORT_STATUS_POWER_SAVE (12)
value PORT_STATUS_TONER_LOW (10)
value PORT_STATUS_TYPE_ERROR (1)
value PORT_STATUS_TYPE_INFO (3)
value PORT_STATUS_TYPE_WARNING (2)
value PORT_STATUS_USER_INTERVENTION (8)
value PORT_STATUS_WARMING_UP (11)
value POSTSCRIPT_DATA (37)
value POSTSCRIPT_IDENTIFY (4117)
value POSTSCRIPT_IGNORE (38)
value POSTSCRIPT_INJECTION (4118)
value POSTSCRIPT_PASSTHROUGH (4115)
value POWERBUTTON_ACTION_INDEX_HIBERNATE (2)
value POWERBUTTON_ACTION_INDEX_NOTHING (0)
value POWERBUTTON_ACTION_INDEX_SHUTDOWN (3)
value POWERBUTTON_ACTION_INDEX_SLEEP (1)
value POWERBUTTON_ACTION_INDEX_TURN_OFF_THE_DISPLAY (4)
value POWERBUTTON_ACTION_VALUE_HIBERNATE (3)
value POWERBUTTON_ACTION_VALUE_NOTHING (0)
value POWERBUTTON_ACTION_VALUE_SHUTDOWN (6)
value POWERBUTTON_ACTION_VALUE_SLEEP (2)
value POWERBUTTON_ACTION_VALUE_TURN_OFF_THE_DISPLAY (8)
value POWER_CONNECTIVITY_IN_STANDBY_DISABLED (0)
value POWER_CONNECTIVITY_IN_STANDBY_ENABLED (1)
value POWER_CONNECTIVITY_IN_STANDBY_SYSTEM_MANAGED (2)
value POWER_DEVICE_IDLE_POLICY_CONSERVATIVE (1)
value POWER_DEVICE_IDLE_POLICY_PERFORMANCE (0)
value POWER_DISCONNECTED_STANDBY_MODE_AGGRESSIVE (1)
value POWER_DISCONNECTED_STANDBY_MODE_NORMAL (0)
value POWER_PLATFORM_ROLE_VERSION (POWER_PLATFORM_ROLE_V2)
value POWER_PLATFORM_ROLE_VERSION_MAX (POWER_PLATFORM_ROLE_V2_MAX)
value POWER_REQUEST_CONTEXT_DETAILED_STRING (DIAGNOSTIC_REASON_DETAILED_STRING)
value POWER_REQUEST_CONTEXT_SIMPLE_STRING (DIAGNOSTIC_REASON_SIMPLE_STRING)
value POWER_REQUEST_CONTEXT_VERSION (DIAGNOSTIC_REASON_VERSION)
value POWER_SYSTEM_MAXIMUM (7)
value PO_THROTTLE_ADAPTIVE (3)
value PO_THROTTLE_CONSTANT (1)
value PO_THROTTLE_DEGRADE (2)
value PO_THROTTLE_MAXIMUM (4)
value PO_THROTTLE_NONE (0)
value PP_ADMIN_PIN (31)
value PP_APPLI_CERT (18)
value PP_CERTCHAIN (9)
value PP_CHANGE_PASSWORD (7)
value PP_CLIENT_HWND (1)
value PP_CONTAINER (6)
value PP_CONTEXT_INFO (11)
value PP_CRYPT_COUNT_KEY_USE (41)
value PP_DELETEKEY (24)
value PP_DISMISS_PIN_UI_SEC (49)
value PP_ENUMALGS (1)
value PP_ENUMALGS_EX (22)
value PP_ENUMCONTAINERS (2)
value PP_ENUMELECTROOTS (26)
value PP_ENUMEX_SIGNING_PROT (40)
value PP_ENUMMANDROOTS (25)
value PP_IMPTYPE (3)
value PP_IS_PFX_EPHEMERAL (50)
value PP_KEYEXCHANGE_ALG (14)
value PP_KEYEXCHANGE_KEYSIZE (12)
value PP_KEYEXCHANGE_PIN (32)
value PP_KEYSET_SEC_DESCR (8)
value PP_KEYSET_TYPE (27)
value PP_KEYSPEC (39)
value PP_KEYSTORAGE (17)
value PP_KEYX_KEYSIZE_INC (35)
value PP_KEY_TYPE_SUBTYPE (10)
value PP_NAME (4)
value PP_PIN_PROMPT_STRING (44)
value PP_PROVTYPE (16)
value PP_ROOT_CERTSTORE (46)
value PP_SECURE_KEYEXCHANGE_PIN (47)
value PP_SECURE_SIGNATURE_PIN (48)
value PP_SESSION_KEYSIZE (20)
value PP_SGC_INFO (37)
value PP_SIGNATURE_ALG (15)
value PP_SIGNATURE_KEYSIZE (13)
value PP_SIGNATURE_PIN (33)
value PP_SIG_KEYSIZE_INC (34)
value PP_SMARTCARD_GUID (45)
value PP_SMARTCARD_READER (43)
value PP_SMARTCARD_READER_ICON (47)
value PP_SYM_KEYSIZE (19)
value PP_UI_PROMPT (21)
value PP_UNIQUE_CONTAINER (36)
value PP_USER_CERTSTORE (42)
value PP_USE_HARDWARE_RNG (38)
value PP_VERSION (5)
value PRAGMA_DEPRECATED_DDK (0)
value PRINTACTION_DOCUMENTDEFAULTS (6)
value PRINTACTION_NETINSTALL (2)
value PRINTACTION_NETINSTALLLINK (3)
value PRINTACTION_OPEN (0)
value PRINTACTION_OPENNETPRN (5)
value PRINTACTION_PROPERTIES (1)
value PRINTACTION_SERVERPROPERTIES (7)
value PRINTACTION_TESTPAGE (4)
value PRINTDLGEXORD (1549)
value PRINTDLGORD (1538)
value PRINTER_CONTROL_PAUSE (1)
value PRINTER_CONTROL_PURGE (3)
value PRINTER_CONTROL_RESUME (2)
value PRINTER_CONTROL_SET_STATUS (4)
value PRINTRATEUNIT_CPS (2)
value PRINTRATEUNIT_IPM (4)
value PRINTRATEUNIT_LPM (3)
value PRINTRATEUNIT_PPM (1)
value PRNSETUPDLGORD (1539)
value PROCESSOR_ARCHITECTURE_ALPHA (2)
value PROCESSOR_ARCHITECTURE_ARM (5)
value PROCESSOR_ARCHITECTURE_INTEL (0)
value PROCESSOR_ARCHITECTURE_MIPS (1)
value PROCESSOR_ARCHITECTURE_MSIL (8)
value PROCESSOR_ARCHITECTURE_NEUTRAL (11)
value PROCESSOR_ARCHITECTURE_PPC (3)
value PROCESSOR_ARCHITECTURE_SHX (4)
value PROCESSOR_DUTY_CYCLING_DISABLED (0)
value PROCESSOR_DUTY_CYCLING_ENABLED (1)
value PROCESSOR_INTEL_PENTIUM (586)
value PROCESSOR_PERF_AUTONOMOUS_MODE_DISABLED (0)
value PROCESSOR_PERF_AUTONOMOUS_MODE_ENABLED (1)
value PROCESSOR_PERF_BOOST_MODE_AGGRESSIVE (2)
value PROCESSOR_PERF_BOOST_MODE_AGGRESSIVE_AT_GUARANTEED (5)
value PROCESSOR_PERF_BOOST_MODE_DISABLED (0)
value PROCESSOR_PERF_BOOST_MODE_EFFICIENT_AGGRESSIVE (4)
value PROCESSOR_PERF_BOOST_MODE_EFFICIENT_AGGRESSIVE_AT_GUARANTEED (6)
value PROCESSOR_PERF_BOOST_MODE_EFFICIENT_ENABLED (3)
value PROCESSOR_PERF_BOOST_MODE_ENABLED (1)
value PROCESSOR_PERF_BOOST_MODE_MAX (PROCESSOR_PERF_BOOST_MODE_EFFICIENT_AGGRESSIVE_AT_GUARANTEED)
value PROCESSOR_PERF_BOOST_POLICY_DISABLED (0)
value PROCESSOR_PERF_BOOST_POLICY_MAX (100)
value PROCESSOR_PERF_ENERGY_PREFERENCE (0)
value PROCESSOR_PERF_MAXIMUM_ACTIVITY_WINDOW (1270000000)
value PROCESSOR_PERF_MINIMUM_ACTIVITY_WINDOW (0)
value PROCESSOR_STRONGARM (2577)
value PROCESSOR_THROTTLE_AUTOMATIC (2)
value PROCESSOR_THROTTLE_DISABLED (0)
value PROCESSOR_THROTTLE_ENABLED (1)
value PROCESS_POWER_THROTTLING_CURRENT_VERSION (1)
value PROC_IDLE_BUCKET_COUNT (6)
value PROC_IDLE_BUCKET_COUNT_EX (16)
value PRODUCT_ID_LENGTH (16)
value PROGRESS_CANCEL (1)
value PROGRESS_CONTINUE (0)
value PROGRESS_QUIET (3)
value PROGRESS_STOP (2)
value PROJFS_PROTOCOL_VERSION (3)
value PROOF_QUALITY (2)
value PROPSHEETHEADER (PROPSHEETHEADERA)
value PROPSHEETPAGE (PROPSHEETPAGEA)
value PROPSHEETPAGE_LATEST (PROPSHEETPAGEA_LATEST)
value PROP_LG_CXDLG (252)
value PROP_LG_CYDLG (218)
value PROP_MED_CXDLG (227)
value PROP_MED_CYDLG (215)
value PROP_SM_CXDLG (212)
value PROP_SM_CYDLG (188)
value PROV_DH_SCHANNEL (18)
value PROV_DSS (3)
value PROV_DSS_DH (13)
value PROV_EC_ECDSA_FULL (16)
value PROV_EC_ECDSA_SIG (14)
value PROV_EC_ECNRA_FULL (17)
value PROV_EC_ECNRA_SIG (15)
value PROV_FORTEZZA (4)
value PROV_INTEL_SEC (22)
value PROV_MS_EXCHANGE (5)
value PROV_REPLACE_OWF (23)
value PROV_RNG (21)
value PROV_RSA_AES (24)
value PROV_RSA_FULL (1)
value PROV_RSA_SCHANNEL (12)
value PROV_RSA_SIG (2)
value PROV_SPYRUS_LYNKS (20)
value PROV_SSL (6)
value PRPC_ENDPOINT_TEMPLATE (PRPC_ENDPOINT_TEMPLATEA)
value PRPC_HTTP_TRANSPORT_CREDENTIALS (PRPC_HTTP_TRANSPORT_CREDENTIALS_A)
value PRPC_INTERFACE_TEMPLATE (PRPC_INTERFACE_TEMPLATEA)
value PSBTN_APPLYNOW (4)
value PSBTN_BACK (0)
value PSBTN_CANCEL (5)
value PSBTN_FINISH (2)
value PSBTN_HELP (6)
value PSBTN_MAX (6)
value PSBTN_NEXT (1)
value PSBTN_OK (3)
value PSCARD_READERSTATE_A (PSCARD_READERSTATEA)
value PSCARD_READERSTATE_W (PSCARD_READERSTATEW)
value PSCB_BUTTONPRESSED (3)
value PSCB_INITIALIZED (1)
value PSCB_PRECREATE (2)
value PSEC_WINNT_AUTH_IDENTITY (PSEC_WINNT_AUTH_IDENTITY_A)
value PSIDENT_GDICENTRIC (0)
value PSIDENT_PSCENTRIC (1)
value PSINJECT_BEGINDEFAULTS (12)
value PSINJECT_BEGINPAGESETUP (101)
value PSINJECT_BEGINPROLOG (14)
value PSINJECT_BEGINSETUP (16)
value PSINJECT_BEGINSTREAM (1)
value PSINJECT_BOUNDINGBOX (9)
value PSINJECT_COMMENTS (11)
value PSINJECT_DOCNEEDEDRES (5)
value PSINJECT_DOCSUPPLIEDRES (6)
value PSINJECT_DOCUMENTPROCESSCOLORS (10)
value PSINJECT_DOCUMENTPROCESSCOLORSATEND (21)
value PSINJECT_ENDDEFAULTS (13)
value PSINJECT_ENDPAGECOMMENTS (107)
value PSINJECT_ENDPAGESETUP (102)
value PSINJECT_ENDPROLOG (15)
value PSINJECT_ENDSETUP (17)
value PSINJECT_ENDSTREAM (20)
value PSINJECT_EOF (19)
value PSINJECT_ORIENTATION (8)
value PSINJECT_PAGEBBOX (106)
value PSINJECT_PAGENUMBER (100)
value PSINJECT_PAGEORDER (7)
value PSINJECT_PAGES (4)
value PSINJECT_PAGESATEND (3)
value PSINJECT_PAGETRAILER (103)
value PSINJECT_PLATECOLOR (104)
value PSINJECT_PSADOBE (2)
value PSINJECT_SHOWPAGE (105)
value PSINJECT_TRAILER (18)
value PSINJECT_VMRESTORE (201)
value PSINJECT_VMSAVE (200)
value PSM_SETBUTTONTEXT (PSM_SETBUTTONTEXTW)
value PSM_SETFINISHTEXT (PSM_SETFINISHTEXTA)
value PSM_SETHEADERSUBTITLE (PSM_SETHEADERSUBTITLEA)
value PSM_SETHEADERTITLE (PSM_SETHEADERTITLEA)
value PSM_SETNEXTTEXT (PSM_SETNEXTTEXTW)
value PSM_SETTITLE (PSM_SETTITLEA)
value PSNRET_INVALID (1)
value PSNRET_INVALID_NOCHANGEPAGE (2)
value PSNRET_MESSAGEHANDLED (3)
value PSNRET_NOERROR (0)
value PSPCB_ADDREF (0)
value PSPCB_CREATE (2)
value PSPCB_RELEASE (1)
value PSPROTOCOL_ASCII (0)
value PSPROTOCOL_BCP (1)
value PSPROTOCOL_BINARY (3)
value PSPROTOCOL_TBCP (2)
value PSWIZB_RESTORE (1)
value PSWIZB_SHOW (0)
value PS_ALTERNATE (8)
value PS_DASH (1)
value PS_DASHDOT (3)
value PS_DASHDOTDOT (4)
value PS_DOT (2)
value PS_INSIDEFRAME (6)
value PS_NULL (5)
value PS_SOLID (0)
value PS_USERSTYLE (7)
value PWR_CRITICALRESUME (3)
value PWR_OK (1)
value PWR_SUSPENDREQUEST (1)
value PWR_SUSPENDRESUME (2)
value QDI_DIBTOSCREEN (4)
value QDI_GETDIBITS (2)
value QDI_SETDIBITS (1)
value QDI_STRETCHDIB (8)
value QOS_GENERAL_ID_BASE (2000)
value QUERYDIBSUPPORT (3073)
value QUERYESCSUPPORT (8)
value QUERYROPSUPPORT (40)
value RANDOM_PADDING (2)
value RASTERCAPS (38)
value RC_BANDING (2)
value RC_BITBLT (1)
value RC_SCALING (4)
value RDH_RECTANGLES (1)
value READ_ATTRIBUTE_BUFFER_SIZE (512)
value READ_THRESHOLD_BUFFER_SIZE (512)
value REASON_LEGACY_API (SHTDN_REASON_LEGACY_API)
value REASON_PLANNED_FLAG (SHTDN_REASON_FLAG_PLANNED)
value REASON_UNKNOWN (SHTDN_REASON_UNKNOWN)
value RECOVERY_DEFAULT_PING_INTERVAL (5000)
value REGISTERWORDENUMPROC (REGISTERWORDENUMPROCA)
value REG_FORCE_UNLOAD (1)
value REG_LATEST_FORMAT (2)
value REG_NO_COMPRESSION (4)
value REG_SECURE_CONNECTION (1)
value REG_STANDARD_FORMAT (1)
value RELATIVE (2)
value REPLACEDLGORD (1541)
value REQUEST_OPLOCK_CURRENT_VERSION (1)
value RESETDEV (7)
value RESTART_MAX_CMD_LINE (1024)
value RESTART_NO_CRASH (1)
value RESTART_NO_HANG (2)
value RESTART_NO_PATCH (4)
value RESTART_NO_REBOOT (8)
value RESTORE_CTM (4100)
value RES_CURSOR (2)
value RES_ICON (1)
value RETRACT_IEPORT (3)
value REVISION_LENGTH (4)
value RGN_AND (1)
value RGN_COPY (5)
value RGN_DIFF (4)
value RGN_ERROR (ERROR)
value RGN_MAX (RGN_COPY)
value RGN_MIN (RGN_AND)
value RGN_OR (2)
value RGN_XOR (3)
value RIM_INPUT (0)
value RIM_INPUTSINK (1)
value RIM_TYPEHID (2)
value RIM_TYPEKEYBOARD (1)
value RIM_TYPEMAX (2)
value RIM_TYPEMOUSE (0)
value RIP_EVENT (9)
value RI_KEY_BREAK (1)
value RI_KEY_MAKE (0)
value RI_KEY_TERMSRV_SET_LED (8)
value ROT_COMPARE_MAX (2048)
value RPCNSAPI (DECLSPEC_IMPORT)
value RPCRTAPI (DECLSPEC_IMPORT)
value RPC_C_AUTHN_CLOUD_AP (36)
value RPC_C_AUTHN_DCE_PRIVATE (1)
value RPC_C_AUTHN_DCE_PUBLIC (2)
value RPC_C_AUTHN_DEC_PUBLIC (4)
value RPC_C_AUTHN_DIGEST (21)
value RPC_C_AUTHN_DPA (17)
value RPC_C_AUTHN_GSS_KERBEROS (16)
value RPC_C_AUTHN_GSS_NEGOTIATE (9)
value RPC_C_AUTHN_GSS_SCHANNEL (14)
value RPC_C_AUTHN_INFO_TYPE_HTTP (1)
value RPC_C_AUTHN_KERNEL (20)
value RPC_C_AUTHN_LEVEL_CALL (3)
value RPC_C_AUTHN_LEVEL_CONNECT (2)
value RPC_C_AUTHN_LEVEL_DEFAULT (0)
value RPC_C_AUTHN_LEVEL_NONE (1)
value RPC_C_AUTHN_LEVEL_PKT (4)
value RPC_C_AUTHN_LEVEL_PKT_INTEGRITY (5)
value RPC_C_AUTHN_LEVEL_PKT_PRIVACY (6)
value RPC_C_AUTHN_LIVEXP_SSP (35)
value RPC_C_AUTHN_LIVE_SSP (32)
value RPC_C_AUTHN_MQ (100)
value RPC_C_AUTHN_MSN (18)
value RPC_C_AUTHN_MSONLINE (82)
value RPC_C_AUTHN_NEGO_EXTENDER (30)
value RPC_C_AUTHN_NONE (0)
value RPC_C_AUTHN_WINNT (10)
value RPC_C_AUTHZ_DCE (2)
value RPC_C_AUTHZ_NAME (1)
value RPC_C_AUTHZ_NONE (0)
value RPC_C_BINDING_DEFAULT_TIMEOUT (5)
value RPC_C_BINDING_INFINITE_TIMEOUT (10)
value RPC_C_BINDING_MAX_TIMEOUT (9)
value RPC_C_BINDING_MIN_TIMEOUT (0)
value RPC_C_BIND_TO_ALL_NICS (1)
value RPC_C_EP_ALL_ELTS (0)
value RPC_C_EP_MATCH_BY_BOTH (3)
value RPC_C_EP_MATCH_BY_IF (1)
value RPC_C_EP_MATCH_BY_OBJ (2)
value RPC_C_HTTP_AUTHN_TARGET_PROXY (2)
value RPC_C_HTTP_AUTHN_TARGET_SERVER (1)
value RPC_C_HTTP_FLAG_ENABLE_CERT_REVOCATION_CHECK (16)
value RPC_C_HTTP_FLAG_IGNORE_CERT_CN_INVALID (8)
value RPC_C_HTTP_FLAG_USE_FIRST_AUTH_SCHEME (2)
value RPC_C_HTTP_FLAG_USE_SSL (1)
value RPC_C_IMP_LEVEL_ANONYMOUS (1)
value RPC_C_IMP_LEVEL_DEFAULT (0)
value RPC_C_IMP_LEVEL_DELEGATE (4)
value RPC_C_IMP_LEVEL_IDENTIFY (2)
value RPC_C_IMP_LEVEL_IMPERSONATE (3)
value RPC_C_INFINITE_TIMEOUT (INFINITE)
value RPC_C_LISTEN_MAX_CALLS_DEFAULT (1234)
value RPC_C_MGMT_INQ_IF_IDS (0)
value RPC_C_MGMT_INQ_PRINC_NAME (1)
value RPC_C_MGMT_INQ_STATS (2)
value RPC_C_MGMT_IS_SERVER_LISTEN (3)
value RPC_C_MGMT_STOP_SERVER_LISTEN (4)
value RPC_C_NS_SYNTAX_DCE (3)
value RPC_C_NS_SYNTAX_DEFAULT (0)
value RPC_C_OPT_ASYNC_BLOCK (15)
value RPC_C_OPT_BINDING_NONCAUSAL (9)
value RPC_C_OPT_CALL_TIMEOUT (12)
value RPC_C_OPT_DONT_LINGER (13)
value RPC_C_OPT_MAX_OPTIONS (17)
value RPC_C_OPT_OPTIMIZE_TIME (16)
value RPC_C_OPT_PRIVATE_BREAK_ON_SUSPEND (3)
value RPC_C_OPT_PRIVATE_DO_NOT_DISTURB (2)
value RPC_C_OPT_PRIVATE_SUPPRESS_WAKE (1)
value RPC_C_OPT_SECURITY_CALLBACK (10)
value RPC_C_OPT_TRANS_SEND_BUFFER_SIZE (5)
value RPC_C_OPT_TRUST_PEER (14)
value RPC_C_OPT_UNIQUE_BINDING (11)
value RPC_C_PARM_BUFFER_LENGTH (2)
value RPC_C_PARM_MAX_PACKET_LENGTH (1)
value RPC_C_PROFILE_ALL_ELT (1)
value RPC_C_PROFILE_ALL_ELTS (RPC_C_PROFILE_ALL_ELT)
value RPC_C_PROFILE_DEFAULT_ELT (0)
value RPC_C_PROFILE_MATCH_BY_BOTH (4)
value RPC_C_PROFILE_MATCH_BY_IF (2)
value RPC_C_PROFILE_MATCH_BY_MBR (3)
value RPC_C_PROTSEQ_MAX_REQS_DEFAULT (10)
value RPC_C_QOS_IDENTITY_DYNAMIC (1)
value RPC_C_QOS_IDENTITY_STATIC (0)
value RPC_C_SECURITY_QOS_VERSION (1L)
value RPC_C_STATS_CALLS_IN (0)
value RPC_C_STATS_CALLS_OUT (1)
value RPC_C_STATS_PKTS_IN (2)
value RPC_C_STATS_PKTS_OUT (3)
value RPC_C_VERS_ALL (1)
value RPC_C_VERS_COMPATIBLE (2)
value RPC_C_VERS_EXACT (3)
value RPC_C_VERS_MAJOR_ONLY (4)
value RPC_C_VERS_UPTO (5)
value RPC_EEINFO_VERSION (1)
value RPC_ENDPOINT_TEMPLATE (RPC_ENDPOINT_TEMPLATEA)
value RPC_HTTP_TRANSPORT_CREDENTIALS (RPC_HTTP_TRANSPORT_CREDENTIALS_A)
value RPC_INTERFACE_TEMPLATE (RPC_INTERFACE_TEMPLATEA)
value RPC_PROTSEQ_VECTOR (RPC_PROTSEQ_VECTORA)
value RPC_PROXY_CONNECTION_TYPE_IN_PROXY (0)
value RPC_PROXY_CONNECTION_TYPE_OUT_PROXY (1)
value RPC_SYSTEM_HANDLE_FREE_ALL (3)
value RPC_SYSTEM_HANDLE_FREE_ERROR_ON_CLOSE (4)
value RPC_SYSTEM_HANDLE_FREE_RETRIEVED (2)
value RPC_SYSTEM_HANDLE_FREE_UNRETRIEVED (1)
value RPC_S_ACCESS_DENIED (ERROR_ACCESS_DENIED)
value RPC_S_ADDRESS_ERROR (1768L)
value RPC_S_ALREADY_LISTENING (1713L)
value RPC_S_ALREADY_REGISTERED (1711L)
value RPC_S_ASYNC_CALL_PENDING (ERROR_IO_PENDING)
value RPC_S_BINDING_HAS_NO_AUTH (1746L)
value RPC_S_BINDING_INCOMPLETE (1819L)
value RPC_S_BUFFER_TOO_SMALL (ERROR_INSUFFICIENT_BUFFER)
value RPC_S_CALL_CANCELLED (1818L)
value RPC_S_CALL_FAILED (1726L)
value RPC_S_CALL_FAILED_DNE (1727L)
value RPC_S_CALL_IN_PROGRESS (1791L)
value RPC_S_CANNOT_SUPPORT (1764L)
value RPC_S_CANT_CREATE_ENDPOINT (1720L)
value RPC_S_COMM_FAILURE (1820L)
value RPC_S_COOKIE_AUTH_FAILED (1833L)
value RPC_S_DO_NOT_DISTURB (1834L)
value RPC_S_DUPLICATE_ENDPOINT (1740L)
value RPC_S_ENTRY_ALREADY_EXISTS (1760L)
value RPC_S_ENTRY_NOT_FOUND (1761L)
value RPC_S_ENTRY_TYPE_MISMATCH (1922L)
value RPC_S_FP_DIV_ZERO (1769L)
value RPC_S_FP_OVERFLOW (1771L)
value RPC_S_FP_UNDERFLOW (1770L)
value RPC_S_GROUP_MEMBER_NOT_FOUND (1898L)
value RPC_S_GRP_ELT_NOT_ADDED (1928L)
value RPC_S_GRP_ELT_NOT_REMOVED (1929L)
value RPC_S_INCOMPLETE_NAME (1755L)
value RPC_S_INTERFACE_NOT_EXPORTED (1924L)
value RPC_S_INTERFACE_NOT_FOUND (1759L)
value RPC_S_INTERNAL_ERROR (1766L)
value RPC_S_INVALID_ARG (ERROR_INVALID_PARAMETER)
value RPC_S_INVALID_ASYNC_CALL (1915L)
value RPC_S_INVALID_ASYNC_HANDLE (1914L)
value RPC_S_INVALID_AUTH_IDENTITY (1749L)
value RPC_S_INVALID_BINDING (1702L)
value RPC_S_INVALID_BOUND (1734L)
value RPC_S_INVALID_ENDPOINT_FORMAT (1706L)
value RPC_S_INVALID_LEVEL (ERROR_INVALID_PARAMETER)
value RPC_S_INVALID_NAF_ID (1763L)
value RPC_S_INVALID_NAME_SYNTAX (1736L)
value RPC_S_INVALID_NETWORK_OPTIONS (1724L)
value RPC_S_INVALID_NET_ADDR (1707L)
value RPC_S_INVALID_OBJECT (1900L)
value RPC_S_INVALID_RPC_PROTSEQ (1704L)
value RPC_S_INVALID_SECURITY_DESC (ERROR_INVALID_SECURITY_DESCR)
value RPC_S_INVALID_STRING_BINDING (1700L)
value RPC_S_INVALID_STRING_UUID (1705L)
value RPC_S_INVALID_TAG (1733L)
value RPC_S_INVALID_TIMEOUT (1709L)
value RPC_S_INVALID_VERS_OPTION (1756L)
value RPC_S_MAX_CALLS_TOO_SMALL (1742L)
value RPC_S_NAME_SERVICE_UNAVAILABLE (1762L)
value RPC_S_NOTHING_TO_EXPORT (1754L)
value RPC_S_NOT_ALL_OBJS_EXPORTED (1923L)
value RPC_S_NOT_ALL_OBJS_UNEXPORTED (1758L)
value RPC_S_NOT_CANCELLED (1826L)
value RPC_S_NOT_ENOUGH_QUOTA (ERROR_NOT_ENOUGH_QUOTA)
value RPC_S_NOT_LISTENING (1715L)
value RPC_S_NOT_RPC_ERROR (1823L)
value RPC_S_NO_BINDINGS (1718L)
value RPC_S_NO_CALL_ACTIVE (1725L)
value RPC_S_NO_CONTEXT_AVAILABLE (1765L)
value RPC_S_NO_ENDPOINT_FOUND (1708L)
value RPC_S_NO_ENTRY_NAME (1735L)
value RPC_S_NO_INTERFACES (1817L)
value RPC_S_NO_MORE_BINDINGS (1806L)
value RPC_S_NO_MORE_MEMBERS (1757L)
value RPC_S_NO_PRINC_NAME (1822L)
value RPC_S_NO_PROTSEQS (1719L)
value RPC_S_NO_PROTSEQS_REGISTERED (1714L)
value RPC_S_OBJECT_NOT_FOUND (1710L)
value RPC_S_OK (ERROR_SUCCESS)
value RPC_S_OUT_OF_MEMORY (ERROR_OUTOFMEMORY)
value RPC_S_OUT_OF_RESOURCES (1721L)
value RPC_S_OUT_OF_THREADS (ERROR_MAX_THRDS_REACHED)
value RPC_S_PRF_ELT_NOT_ADDED (1926L)
value RPC_S_PRF_ELT_NOT_REMOVED (1927L)
value RPC_S_PROCNUM_OUT_OF_RANGE (1745L)
value RPC_S_PROFILE_NOT_ADDED (1925L)
value RPC_S_PROTOCOL_ERROR (1728L)
value RPC_S_PROTSEQ_NOT_FOUND (1744L)
value RPC_S_PROTSEQ_NOT_SUPPORTED (1703L)
value RPC_S_PROXY_ACCESS_DENIED (1729L)
value RPC_S_RUNTIME_UNINITIALIZED (ERROR_INVALID_FUNCTION)
value RPC_S_SEC_PKG_ERROR (1825L)
value RPC_S_SEND_INCOMPLETE (1913L)
value RPC_S_SERVER_OUT_OF_MEMORY (ERROR_NOT_ENOUGH_SERVER_MEMORY)
value RPC_S_SERVER_TOO_BUSY (1723L)
value RPC_S_SERVER_UNAVAILABLE (1722L)
value RPC_S_STRING_TOO_LONG (1743L)
value RPC_S_SYSTEM_HANDLE_COUNT_EXCEEDED (1835L)
value RPC_S_SYSTEM_HANDLE_TYPE_MISMATCH (1836L)
value RPC_S_TIMEOUT (ERROR_TIMEOUT)
value RPC_S_TYPE_ALREADY_REGISTERED (1712L)
value RPC_S_UNKNOWN_AUTHN_LEVEL (1748L)
value RPC_S_UNKNOWN_AUTHN_SERVICE (1747L)
value RPC_S_UNKNOWN_AUTHN_TYPE (1741L)
value RPC_S_UNKNOWN_AUTHZ_SERVICE (1750L)
value RPC_S_UNKNOWN_IF (1717L)
value RPC_S_UNKNOWN_MGR_TYPE (1716L)
value RPC_S_UNKNOWN_PRINCIPAL (ERROR_NONE_MAPPED)
value RPC_S_UNSUPPORTED_AUTHN_LEVEL (1821L)
value RPC_S_UNSUPPORTED_NAME_SYNTAX (1737L)
value RPC_S_UNSUPPORTED_TRANS_SYN (1730L)
value RPC_S_UNSUPPORTED_TYPE (1732L)
value RPC_S_UUID_LOCAL_ONLY (1824L)
value RPC_S_UUID_NO_ADDRESS (1739L)
value RPC_S_WRONG_KIND_OF_BINDING (1701L)
value RPC_S_ZERO_DIVIDE (1767L)
value RPC_X_BAD_STUB_DATA (1783L)
value RPC_X_BYTE_COUNT_TOO_SMALL (1782L)
value RPC_X_ENUM_VALUE_OUT_OF_RANGE (1781L)
value RPC_X_ENUM_VALUE_TOO_LARGE (RPC_X_ENUM_VALUE_OUT_OF_RANGE)
value RPC_X_INVALID_BOUND (RPC_S_INVALID_BOUND)
value RPC_X_INVALID_BUFFER (ERROR_INVALID_USER_BUFFER)
value RPC_X_INVALID_ES_ACTION (1827L)
value RPC_X_INVALID_PIPE_OBJECT (1830L)
value RPC_X_INVALID_PIPE_OPERATION (RPC_X_WRONG_PIPE_ORDER)
value RPC_X_INVALID_TAG (RPC_S_INVALID_TAG)
value RPC_X_NO_MEMORY (RPC_S_OUT_OF_MEMORY)
value RPC_X_NO_MORE_ENTRIES (1772L)
value RPC_X_NULL_REF_POINTER (1780L)
value RPC_X_PIPE_APP_MEMORY (ERROR_OUTOFMEMORY)
value RPC_X_PIPE_CLOSED (1916L)
value RPC_X_PIPE_DISCIPLINE_ERROR (1917L)
value RPC_X_PIPE_EMPTY (1918L)
value RPC_X_SS_CANNOT_GET_CALL_HANDLE (1779L)
value RPC_X_SS_CHAR_TRANS_OPEN_FAIL (1773L)
value RPC_X_SS_CHAR_TRANS_SHORT_FILE (1774L)
value RPC_X_SS_CONTEXT_DAMAGED (1777L)
value RPC_X_SS_CONTEXT_MISMATCH (ERROR_INVALID_HANDLE)
value RPC_X_SS_HANDLES_MISMATCH (1778L)
value RPC_X_SS_IN_NULL_CONTEXT (1775L)
value RPC_X_WRONG_ES_VERSION (1828L)
value RPC_X_WRONG_PIPE_ORDER (1831L)
value RPC_X_WRONG_PIPE_VERSION (1832L)
value RPC_X_WRONG_STUB_VERSION (1829L)
value RTL_CORRELATION_VECTOR_STRING_LENGTH (129)
value RTL_CORRELATION_VECTOR_VERSION_CURRENT (RTL_CORRELATION_VECTOR_VERSION_2)
value RTL_RUN_ONCE_CTX_RESERVED_BITS (2)
value RUNDLGORD (1545)
value RUSSIAN_CHARSET (204)
value SAVE_CTM (4101)
value SB_BOTH (3)
value SB_BOTTOM (7)
value SB_CTL (2)
value SB_ENDSCROLL (8)
value SB_HORZ (0)
value SB_LEFT (6)
value SB_LINEDOWN (1)
value SB_LINELEFT (0)
value SB_LINERIGHT (1)
value SB_LINEUP (0)
value SB_PAGEDOWN (3)
value SB_PAGELEFT (2)
value SB_PAGERIGHT (3)
value SB_PAGEUP (2)
value SB_RIGHT (7)
value SB_THUMBPOSITION (4)
value SB_THUMBTRACK (5)
value SB_TOP (6)
value SB_VERT (1)
value SCALINGFACTORX (114)
value SCALINGFACTORY (115)
value SCARD_ABSENT (1)
value SCARD_ATR_LENGTH (33)
value SCARD_ATTR_DEVICE_FRIENDLY_NAME (SCARD_ATTR_DEVICE_FRIENDLY_NAME_A)
value SCARD_ATTR_DEVICE_SYSTEM_NAME (SCARD_ATTR_DEVICE_SYSTEM_NAME_A)
value SCARD_CLASS_COMMUNICATIONS (2)
value SCARD_CLASS_ICC_STATE (9)
value SCARD_CLASS_IFD_PROTOCOL (8)
value SCARD_CLASS_MECHANICAL (6)
value SCARD_CLASS_POWER_MGMT (4)
value SCARD_CLASS_PROTOCOL (3)
value SCARD_CLASS_SECURITY (5)
value SCARD_CLASS_VENDOR_DEFINED (7)
value SCARD_CLASS_VENDOR_INFO (1)
value SCARD_COLD_RESET (1)
value SCARD_EJECT_CARD (3)
value SCARD_LEAVE_CARD (0)
value SCARD_NEGOTIABLE (5)
value SCARD_POWERED (4)
value SCARD_POWER_DOWN (0)
value SCARD_PRESENT (2)
value SCARD_PROVIDER_CSP (2)
value SCARD_PROVIDER_KSP (3)
value SCARD_PROVIDER_PRIMARY (1)
value SCARD_READERSTATE_A (SCARD_READERSTATEA)
value SCARD_READERSTATE_W (SCARD_READERSTATEW)
value SCARD_RESET_CARD (1)
value SCARD_SCOPE_SYSTEM (2)
value SCARD_SCOPE_TERMINAL (1)
value SCARD_SCOPE_USER (0)
value SCARD_SHARE_DIRECT (3)
value SCARD_SHARE_EXCLUSIVE (1)
value SCARD_SHARE_SHARED (2)
value SCARD_SPECIFIC (6)
value SCARD_SWALLOWED (3)
value SCARD_S_SUCCESS (NO_ERROR)
value SCARD_UNKNOWN (0)
value SCARD_UNPOWER_CARD (2)
value SCARD_WARM_RESET (2)
value SCHAR_MAX (127)
value SCHED_E_SERVICE_NOT_LOCALSYSTEM (6200L)
value SCM_MAX_SYMLINK_LEN_IN_CHARS (256)
value SCM_PD_FIRMWARE_REVISION_LENGTH_BYTES (32)
value SCM_PD_MAX_OPERATIONAL_STATUS (16)
value SCM_PD_MEMORY_SIZE_UNKNOWN (MAXDWORD64)
value SCM_PD_PROPERTY_NAME_LENGTH_IN_CHARS (128)
value SCM_REGION_SPA_UNKNOWN (MAXDWORD64)
value SCS_DOS_BINARY (1)
value SCS_PIF_BINARY (3)
value SCS_POSIX_BINARY (4)
value SCS_THIS_PLATFORM_BINARY (SCS_64BIT_BINARY)
value SCS_WOW_BINARY (2)
value SC_GROUP_IDENTIFIER (SC_GROUP_IDENTIFIERA)
value SC_ICON (SC_MINIMIZE)
value SC_ZOOM (SC_MAXIMIZE)
value SD_GLOBAL_CHANGE_TYPE_MACHINE_SID (1)
value SECURITY_MANDATORY_MAXIMUM_USER_RID (SECURITY_MANDATORY_SYSTEM_RID)
value SECURITY_SERVER_LOGON_RID (SECURITY_ENTERPRISE_CONTROLLERS_RID)
value SEC_E_NOT_SUPPORTED (SEC_E_UNSUPPORTED_FUNCTION)
value SEC_E_NO_SPM (SEC_E_INTERNAL_ERROR)
value SEC_WINNT_AUTH_IDENTITY (SEC_WINNT_AUTH_IDENTITY_A)
value SEEK_CUR (1)
value SEEK_END (2)
value SEEK_SET (0)
value SEE_MASK_FLAG_DDEWAIT (SEE_MASK_NOASYNC)
value SELECTDIB (41)
value SELECTPAPERSOURCE (18)
value SERIAL_NUMBER_LENGTH (32)
value SERVICES_ACTIVE_DATABASE (SERVICES_ACTIVE_DATABASEA)
value SERVICES_FAILED_DATABASE (SERVICES_FAILED_DATABASEA)
value SERVICE_CONFIG_DELAYED_AUTO_START_INFO (3)
value SERVICE_CONFIG_DESCRIPTION (1)
value SERVICE_CONFIG_FAILURE_ACTIONS (2)
value SERVICE_CONFIG_FAILURE_ACTIONS_FLAG (4)
value SERVICE_CONFIG_LAUNCH_PROTECTED (12)
value SERVICE_CONFIG_PREFERRED_NODE (9)
value SERVICE_CONFIG_PRESHUTDOWN_INFO (7)
value SERVICE_CONFIG_REQUIRED_PRIVILEGES_INFO (6)
value SERVICE_CONFIG_SERVICE_SID_INFO (5)
value SERVICE_CONFIG_TRIGGER_INFO (8)
value SERVICE_CONTROL_STATUS_REASON_INFO (1)
value SERVICE_DYNAMIC_INFORMATION_LEVEL_START_REASON (1)
value SERVICE_LAUNCH_PROTECTED_ANTIMALWARE_LIGHT (3)
value SERVICE_LAUNCH_PROTECTED_NONE (0)
value SERVICE_LAUNCH_PROTECTED_WINDOWS (1)
value SERVICE_LAUNCH_PROTECTED_WINDOWS_LIGHT (2)
value SERVICE_MAIN_FUNCTION (SERVICE_MAIN_FUNCTIONA)
value SERVICE_NOTIFY_STATUS_CHANGE (SERVICE_NOTIFY_STATUS_CHANGE_2)
value SERVICE_TRIGGER_ACTION_SERVICE_START (1)
value SERVICE_TRIGGER_ACTION_SERVICE_STOP (2)
value SERVICE_TRIGGER_DATA_TYPE_BINARY (1)
value SERVICE_TRIGGER_DATA_TYPE_KEYWORD_ALL (5)
value SERVICE_TRIGGER_DATA_TYPE_KEYWORD_ANY (4)
value SERVICE_TRIGGER_DATA_TYPE_LEVEL (3)
value SERVICE_TRIGGER_DATA_TYPE_STRING (2)
value SERVICE_TRIGGER_TYPE_AGGREGATE (30)
value SERVICE_TRIGGER_TYPE_CUSTOM (20)
value SERVICE_TRIGGER_TYPE_CUSTOM_SYSTEM_STATE_CHANGE (7)
value SERVICE_TRIGGER_TYPE_DEVICE_INTERFACE_ARRIVAL (1)
value SERVICE_TRIGGER_TYPE_DOMAIN_JOIN (3)
value SERVICE_TRIGGER_TYPE_FIREWALL_PORT_EVENT (4)
value SERVICE_TRIGGER_TYPE_GROUP_POLICY (5)
value SERVICE_TRIGGER_TYPE_IP_ADDRESS_AVAILABILITY (2)
value SERVICE_TRIGGER_TYPE_NETWORK_ENDPOINT (6)
value SERVICE_TYPE_VALUE_OBJECTID (SERVICE_TYPE_VALUE_OBJECTIDA)
value SERVICE_TYPE_VALUE_SAPID (SERVICE_TYPE_VALUE_SAPIDA)
value SERVICE_TYPE_VALUE_TCPPORT (SERVICE_TYPE_VALUE_TCPPORTA)
value SERVICE_TYPE_VALUE_UDPPORT (SERVICE_TYPE_VALUE_UDPPORTA)
value SETABORTPROC (9)
value SETALLJUSTVALUES (771)
value SETBREAK (8)
value SETCHARSET (772)
value SETCOLORTABLE (4)
value SETCOPYCOUNT (17)
value SETDIBSCALING (32)
value SETDTR (5)
value SETKERNTRACK (770)
value SETLINECAP (21)
value SETLINEJOIN (22)
value SETMITERLIMIT (23)
value SETRGBSTRING (SETRGBSTRINGA)
value SETRTS (3)
value SETXOFF (1)
value SETXON (2)
value SET_ARC_DIRECTION (4102)
value SET_BACKGROUND_COLOR (4103)
value SET_BOUNDS (4109)
value SET_CLIP_BOX (4108)
value SET_MIRROR_MODE (4110)
value SET_POLY_MODE (4104)
value SET_SCREEN_ANGLE (4105)
value SET_SPREAD (4106)
value SET_TAPE_DRIVE_INFORMATION (1)
value SET_TAPE_MEDIA_INFORMATION (0)
value SEVERITY_ERROR (1)
value SEVERITY_SUCCESS (0)
value SE_ERR_ACCESSDENIED (5)
value SE_ERR_ASSOCINCOMPLETE (27)
value SE_ERR_DDEBUSY (30)
value SE_ERR_DDEFAIL (29)
value SE_ERR_DDETIMEOUT (28)
value SE_ERR_DLLNOTFOUND (32)
value SE_ERR_FNF (2)
value SE_ERR_NOASSOC (31)
value SE_ERR_OOM (8)
value SE_ERR_PNF (3)
value SE_ERR_SHARE (26)
value SE_SIGNING_LEVEL_ANTIMALWARE (SE_SIGNING_LEVEL_CUSTOM_3)
value SE_SIGNING_LEVEL_DEVELOPER (SE_SIGNING_LEVEL_CUSTOM_1)
value SHADEBLENDCAPS (120)
value SHAREVISTRING (SHAREVISTRINGA)
value SHGSI_ICON (SHGFI_ICON)
value SHGSI_ICONLOCATION (0)
value SHGSI_LARGEICON (SHGFI_LARGEICON)
value SHGSI_LINKOVERLAY (SHGFI_LINKOVERLAY)
value SHGSI_SELECTED (SHGFI_SELECTED)
value SHGSI_SHELLICONSIZE (SHGFI_SHELLICONSIZE)
value SHGSI_SMALLICON (SHGFI_SMALLICON)
value SHGSI_SYSICONINDEX (SHGFI_SYSICONINDEX)
value SHIFTJIS_CHARSET (128)
value SHIL_EXTRALARGE (2)
value SHIL_JUMBO (4)
value SHIL_LARGE (0)
value SHIL_LAST (SHIL_JUMBO)
value SHIL_SMALL (1)
value SHIL_SYSSMALL (3)
value SHOW_FULLSCREEN (3)
value SHOW_ICONWINDOW (2)
value SHOW_OPENNOACTIVATE (4)
value SHOW_OPENWINDOW (1)
value SHRT_MAX (32767)
value SHTDN_REASON_UNKNOWN (SHTDN_REASON_MINOR_NONE)
value SHUTDOWN_TYPE_LEN (32)
value SID_HASH_SIZE (32)
value SIMPLEREGION (2)
value SIZEFULLSCREEN (SIZE_MAXIMIZED)
value SIZEICONIC (SIZE_MINIMIZED)
value SIZENORMAL (SIZE_RESTORED)
value SIZEOF_RFPO_DATA (16)
value SIZEPALETTE (104)
value SIZEZOOMHIDE (SIZE_MAXHIDE)
value SIZEZOOMSHOW (SIZE_MAXSHOW)
value SIZE_MAXHIDE (4)
value SIZE_MAXIMIZED (2)
value SIZE_MAXSHOW (3)
value SIZE_MINIMIZED (1)
value SIZE_RESTORED (0)
value SMART_ABORT_OFFLINE_SELFTEST (127)
value SMART_ERROR_NO_MEM (7)
value SMART_EXTENDED_SELFTEST_CAPTIVE (130)
value SMART_EXTENDED_SELFTEST_OFFLINE (2)
value SMART_IDE_ERROR (1)
value SMART_INVALID_BUFFER (4)
value SMART_INVALID_COMMAND (3)
value SMART_INVALID_DRIVE (5)
value SMART_INVALID_FLAG (2)
value SMART_INVALID_IOCTL (6)
value SMART_INVALID_REGISTER (8)
value SMART_LOG_SECTOR_SIZE (512)
value SMART_NOT_SUPPORTED (9)
value SMART_NO_ERROR (0)
value SMART_NO_IDE_DEVICE (10)
value SMART_OFFLINE_ROUTINE_OFFLINE (0)
value SMART_SHORT_SELFTEST_CAPTIVE (129)
value SMART_SHORT_SELFTEST_OFFLINE (1)
value SMT_UNPARKING_POLICY_CORE (0)
value SMT_UNPARKING_POLICY_CORE_PER_THREAD (1)
value SMT_UNPARKING_POLICY_LP_ROUNDROBIN (2)
value SMT_UNPARKING_POLICY_LP_SEQUENTIAL (3)
value SM_ARRANGE (56)
value SM_CLEANBOOT (67)
value SM_CMETRICS (97)
value SM_CMONITORS (80)
value SM_CMOUSEBUTTONS (43)
value SM_CXBORDER (5)
value SM_CXCURSOR (13)
value SM_CXDLGFRAME (7)
value SM_CXDOUBLECLK (36)
value SM_CXDRAG (68)
value SM_CXEDGE (45)
value SM_CXFIXEDFRAME (SM_CXDLGFRAME)
value SM_CXFOCUSBORDER (83)
value SM_CXFRAME (32)
value SM_CXFULLSCREEN (16)
value SM_CXHSCROLL (21)
value SM_CXHTHUMB (10)
value SM_CXICON (11)
value SM_CXICONSPACING (38)
value SM_CXMAXIMIZED (61)
value SM_CXMAXTRACK (59)
value SM_CXMENUCHECK (71)
value SM_CXMENUSIZE (54)
value SM_CXMIN (28)
value SM_CXMINIMIZED (57)
value SM_CXMINSPACING (47)
value SM_CXMINTRACK (34)
value SM_CXPADDEDBORDER (92)
value SM_CXSCREEN (0)
value SM_CXSIZE (30)
value SM_CXSIZEFRAME (SM_CXFRAME)
value SM_CXSMICON (49)
value SM_CXSMSIZE (52)
value SM_CXVIRTUALSCREEN (78)
value SM_CXVSCROLL (2)
value SM_CYBORDER (6)
value SM_CYCAPTION (4)
value SM_CYCURSOR (14)
value SM_CYDLGFRAME (8)
value SM_CYDOUBLECLK (37)
value SM_CYDRAG (69)
value SM_CYEDGE (46)
value SM_CYFIXEDFRAME (SM_CYDLGFRAME)
value SM_CYFOCUSBORDER (84)
value SM_CYFRAME (33)
value SM_CYFULLSCREEN (17)
value SM_CYHSCROLL (3)
value SM_CYICON (12)
value SM_CYICONSPACING (39)
value SM_CYKANJIWINDOW (18)
value SM_CYMAXIMIZED (62)
value SM_CYMAXTRACK (60)
value SM_CYMENU (15)
value SM_CYMENUCHECK (72)
value SM_CYMENUSIZE (55)
value SM_CYMIN (29)
value SM_CYMINIMIZED (58)
value SM_CYMINSPACING (48)
value SM_CYMINTRACK (35)
value SM_CYSCREEN (1)
value SM_CYSIZE (31)
value SM_CYSIZEFRAME (SM_CYFRAME)
value SM_CYSMCAPTION (51)
value SM_CYSMICON (50)
value SM_CYSMSIZE (53)
value SM_CYVIRTUALSCREEN (79)
value SM_CYVSCROLL (20)
value SM_CYVTHUMB (9)
value SM_DBCSENABLED (42)
value SM_DEBUG (22)
value SM_DIGITIZER (94)
value SM_IMMENABLED (82)
value SM_MAXIMUMTOUCHES (95)
value SM_MEDIACENTER (87)
value SM_MENUDROPALIGNMENT (40)
value SM_MIDEASTENABLED (74)
value SM_MOUSEHORIZONTALWHEELPRESENT (91)
value SM_MOUSEPRESENT (19)
value SM_MOUSEWHEELPRESENT (75)
value SM_NETWORK (63)
value SM_PENWINDOWS (41)
value SM_SAMEDISPLAYFORMAT (81)
value SM_SECURE (44)
value SM_SHOWSOUNDS (70)
value SM_SLOWMACHINE (73)
value SM_STARTER (88)
value SM_SWAPBUTTON (23)
value SM_TABLETPC (86)
value SM_XVIRTUALSCREEN (76)
value SM_YVIRTUALSCREEN (77)
value SNAPSHOT_POLICY_ALWAYS (1)
value SNAPSHOT_POLICY_NEVER (0)
value SNAPSHOT_POLICY_UNPLANNED (2)
value SND_ALIAS_START (0)
value SOCK_DGRAM (2)
value SOCK_NOTIFY_EVENT_HANGUP (SOCK_NOTIFY_REGISTER_EVENT_HANGUP)
value SOCK_NOTIFY_EVENT_IN (SOCK_NOTIFY_REGISTER_EVENT_IN)
value SOCK_NOTIFY_EVENT_OUT (SOCK_NOTIFY_REGISTER_EVENT_OUT)
value SOCK_RAW (3)
value SOCK_RDM (4)
value SOCK_SEQPACKET (5)
value SOCK_STREAM (1)
value SOUND_SYSTEM_APPEND (14)
value SOUND_SYSTEM_APPSTART (12)
value SOUND_SYSTEM_BEEP (3)
value SOUND_SYSTEM_ERROR (4)
value SOUND_SYSTEM_FAULT (13)
value SOUND_SYSTEM_INFORMATION (7)
value SOUND_SYSTEM_MAXIMIZE (8)
value SOUND_SYSTEM_MENUCOMMAND (15)
value SOUND_SYSTEM_MENUPOPUP (16)
value SOUND_SYSTEM_MINIMIZE (9)
value SOUND_SYSTEM_QUESTION (5)
value SOUND_SYSTEM_RESTOREDOWN (11)
value SOUND_SYSTEM_RESTOREUP (10)
value SOUND_SYSTEM_SHUTDOWN (2)
value SOUND_SYSTEM_STARTUP (1)
value SOUND_SYSTEM_WARNING (6)
value SO_PROTOCOL_INFO (SO_PROTOCOL_INFOA)
value SPACEPARITY (4)
value SPIF_SENDCHANGE (SPIF_SENDWININICHANGE)
value SPI_GETMENUUNDERLINES (SPI_GETKEYBOARDCUES)
value SPI_SCREENSAVERRUNNING (SPI_SETSCREENSAVERRUNNING)
value SPI_SETMENUUNDERLINES (SPI_SETKEYBOARDCUES)
value SRB_TYPE_SCSI_REQUEST_BLOCK (0)
value SRB_TYPE_STORAGE_REQUEST_BLOCK (1)
value SRWLOCK_INIT (RTL_SRWLOCK_INIT)
value SSGF_DISPLAY (3)
value SSGF_NONE (0)
value SSL_HPKP_HEADER_COUNT (2)
value SSL_HPKP_PKP_HEADER_INDEX (0)
value SSL_HPKP_PKP_RO_HEADER_INDEX (1)
value SSL_KEY_PIN_ERROR_TEXT_LENGTH (512)
value SSTF_BORDER (2)
value SSTF_CHARS (1)
value SSTF_DISPLAY (3)
value SSTF_NONE (0)
value SSWF_CUSTOM (4)
value SSWF_DISPLAY (3)
value SSWF_NONE (0)
value SSWF_TITLE (1)
value SSWF_WINDOW (2)
value STARTDOC (10)
value STATE_SYSTEM_INDETERMINATE (STATE_SYSTEM_MIXED)
value STGFMT_ANY (4)
value STGFMT_DOCFILE (5)
value STGFMT_DOCUMENT (0)
value STGFMT_FILE (3)
value STGFMT_NATIVE (1)
value STGFMT_STORAGE (0)
value STGOPTIONS_VERSION (2)
value STILL_ACTIVE (STATUS_PENDING)
value STKFORCEINLINE (FORCEINLINE)
value STN_CLICKED (0)
value STN_DBLCLK (1)
value STN_DISABLE (3)
value STN_ENABLE (2)
value STOCK_LAST (19)
value STORAGE_DEVICE_MAX_OPERATIONAL_STATUS (16)
value STORAGE_DEVICE_NUMA_NODE_UNKNOWN (MAXDWORD)
value STORAGE_HW_FIRMWARE_REVISION_LENGTH (16)
value STORAGE_OFFLOAD_MAX_TOKEN_LENGTH (512)
value STORAGE_RPMB_MINIMUM_RELIABLE_WRITE_SIZE (512)
value STORATTRIBUTE_MANAGEMENT_STATE (1)
value STORATTRIBUTE_NONE (0)
value STORE_ERROR_LICENSE_REVOKED (15864L)
value STORE_ERROR_PENDING_COM_TRANSACTION (15863L)
value STORE_ERROR_UNLICENSED (15861L)
value STORE_ERROR_UNLICENSED_USER (15862L)
value STRETCHBLT (2048)
value STRETCH_ANDSCANS (BLACKONWHITE)
value STRETCH_DELETESCANS (COLORONCOLOR)
value STRETCH_HALFTONE (HALFTONE)
value STRETCH_ORSCANS (WHITEONBLACK)
value STRICT (1)
value STRUNCATE (80)
value STYLE_DESCRIPTION_SIZE (32)
value SUPPORT_LANG_NUMBER (32)
value SWP_DRAWFRAME (SWP_FRAMECHANGED)
value SWP_NOREPOSITION (SWP_NOOWNERZORDER)
value SW_FORCEMINIMIZE (11)
value SW_HIDE (0)
value SW_MAX (11)
value SW_MAXIMIZE (3)
value SW_MINIMIZE (6)
value SW_NORMAL (1)
value SW_OTHERUNZOOM (4)
value SW_OTHERZOOM (2)
value SW_PARENTCLOSING (1)
value SW_PARENTOPENING (3)
value SW_RESTORE (9)
value SW_SHOW (5)
value SW_SHOWDEFAULT (10)
value SW_SHOWMAXIMIZED (3)
value SW_SHOWMINIMIZED (2)
value SW_SHOWMINNOACTIVE (7)
value SW_SHOWNA (8)
value SW_SHOWNOACTIVATE (4)
value SW_SHOWNORMAL (1)
value SYMBOL_CHARSET (2)
value SYSPAL_ERROR (0)
value SYSPAL_NOSTATIC (2)
value SYSPAL_STATIC (1)
value SYSRGN (4)
value SYSTEM_CACHE_ALIGNMENT_SIZE (X86_CACHE_ALIGNMENT_SIZE)
value SYSTEM_FIXED_FONT (16)
value SYSTEM_FONT (13)
value SYS_OPEN (_SYS_OPEN)
value S_ALLTHRESHOLD (2)
value S_ASYNCHRONOUS (MK_S_ASYNCHRONOUS)
value S_IEXEC (_S_IEXEC)
value S_IFCHR (_S_IFCHR)
value S_IFDIR (_S_IFDIR)
value S_IFMT (_S_IFMT)
value S_IFREG (_S_IFREG)
value S_IREAD (_S_IREAD)
value S_IWRITE (_S_IWRITE)
value S_LEGATO (1)
value S_NORMAL (0)
value S_PERIODVOICE (3)
value S_QUEUEEMPTY (0)
value S_STACCATO (2)
value S_THRESHOLD (1)
value S_WHITEVOICE (7)
value TAPE_ABSOLUTE_BLOCK (1L)
value TAPE_ABSOLUTE_POSITION (0cL)
value TAPE_CHECK_FOR_DRIVE_PROBLEM (2L)
value TAPE_ERASE_LONG (1L)
value TAPE_ERASE_SHORT (0cL)
value TAPE_FILEMARKS (1L)
value TAPE_FIXED_PARTITIONS (0cL)
value TAPE_FORMAT (5L)
value TAPE_INITIATOR_PARTITIONS (2L)
value TAPE_LOAD (0cL)
value TAPE_LOCK (3L)
value TAPE_LOGICAL_BLOCK (2L)
value TAPE_LOGICAL_POSITION (1L)
value TAPE_LONG_FILEMARKS (3L)
value TAPE_PSEUDO_LOGICAL_BLOCK (3L)
value TAPE_PSEUDO_LOGICAL_POSITION (2L)
value TAPE_QUERY_DEVICE_ERROR_DATA (4L)
value TAPE_QUERY_DRIVE_PARAMETERS (0cL)
value TAPE_QUERY_IO_ERROR_DATA (3L)
value TAPE_QUERY_MEDIA_CAPACITY (1L)
value TAPE_RESET_STATISTICS (2L)
value TAPE_RETURN_ENV_INFO (1L)
value TAPE_RETURN_STATISTICS (0cL)
value TAPE_REWIND (0cL)
value TAPE_SELECT_PARTITIONS (1L)
value TAPE_SETMARKS (0cL)
value TAPE_SHORT_FILEMARKS (2L)
value TAPE_SPACE_END_OF_DATA (4L)
value TAPE_SPACE_FILEMARKS (6L)
value TAPE_SPACE_RELATIVE_BLOCKS (5L)
value TAPE_SPACE_SEQUENTIAL_FMKS (7L)
value TAPE_SPACE_SEQUENTIAL_SMKS (9L)
value TAPE_SPACE_SETMARKS (8L)
value TAPE_TENSION (2L)
value TAPE_UNLOAD (1L)
value TAPE_UNLOCK (4L)
value TA_BASELINE (24)
value TA_BOTTOM (8)
value TA_CENTER (6)
value TA_LEFT (0)
value TA_NOUPDATECP (0)
value TA_RIGHT (2)
value TA_RTLREADING (256)
value TA_TOP (0)
value TA_UPDATECP (1)
value TCI_SRCCHARSET (1)
value TCI_SRCCODEPAGE (2)
value TCI_SRCFONTSIG (3)
value TC_DEVICEDUMP_SUBSECTION_DESC_LENGTH (16)
value TC_GP_TRAP (2)
value TC_HARDERR (1)
value TC_NONCONF_BORROW (0)
value TC_NONCONF_BORROW_PLUS (3)
value TC_NONCONF_DISCARD (2)
value TC_NONCONF_SHAPE (1)
value TC_NORMAL (0)
value TC_PUBLIC_DEVICEDUMP_CONTENT_GPLOG_MAX (16)
value TC_SIGNAL (3)
value TECHNOLOGY (2)
value TELEMETRY_COMMAND_SIZE (16)
value TEXTCAPS (34)
value THAI_CHARSET (222)
value THREAD_BASE_PRIORITY_LOWRT (15)
value THREAD_BASE_PRIORITY_MAX (2)
value THREAD_DYNAMIC_CODE_ALLOW (1)
value THREAD_POWER_THROTTLING_CURRENT_VERSION (1)
value THREAD_PRIORITY_HIGHEST (THREAD_BASE_PRIORITY_MAX)
value THREAD_PRIORITY_IDLE (THREAD_BASE_PRIORITY_IDLE)
value THREAD_PRIORITY_LOWEST (THREAD_BASE_PRIORITY_MIN)
value THREAD_PRIORITY_NORMAL (0)
value THREAD_PRIORITY_TIME_CRITICAL (THREAD_BASE_PRIORITY_LOWRT)
value TIMEFMT_ENUMPROC (TIMEFMT_ENUMPROCA)
value TIMERR_BASE (96)
value TIMESTAMP_FAILURE_BAD_ALG (0)
value TIMESTAMP_FAILURE_BAD_FORMAT (5)
value TIMESTAMP_FAILURE_BAD_REQUEST (2)
value TIMESTAMP_FAILURE_EXTENSION_NOT_SUPPORTED (16)
value TIMESTAMP_FAILURE_INFO_NOT_AVAILABLE (17)
value TIMESTAMP_FAILURE_POLICY_NOT_SUPPORTED (15)
value TIMESTAMP_FAILURE_SYSTEM_FAILURE (25)
value TIMESTAMP_FAILURE_TIME_NOT_AVAILABLE (14)
value TIMESTAMP_STATUS_GRANTED (0)
value TIMESTAMP_STATUS_GRANTED_WITH_MODS (1)
value TIMESTAMP_STATUS_REJECTED (2)
value TIMESTAMP_STATUS_REVOCATION_WARNING (4)
value TIMESTAMP_STATUS_REVOKED (5)
value TIMESTAMP_STATUS_WAITING (3)
value TIMESTAMP_VERSION (1)
value TIME_UTC (1)
value TIME_ZONE_ID_DAYLIGHT (2)
value TIME_ZONE_ID_STANDARD (1)
value TIME_ZONE_ID_UNKNOWN (0)
value TLS_MINIMUM_AVAILABLE (64)
value TMP_MAX (_CRT_INT_MAX)
value TMP_MAX_S (TMP_MAX)
value TOKEN_ACCESS_PSEUDO_HANDLE (TOKEN_ACCESS_PSEUDO_HANDLE_WIN8)
value TOKEN_SOURCE_LENGTH (8)
value TOUCHPREDICTIONPARAMETERS_DEFAULT_LATENCY (8)
value TOUCHPREDICTIONPARAMETERS_DEFAULT_SAMPLETIME (8)
value TOUCHPREDICTIONPARAMETERS_DEFAULT_USE_HW_TIMESTAMP (1)
value TRANSFORM_CTM (4107)
value TRANSPARENT (1)
value TRUE (1)
value TRUNCATE_EXISTING (5)
value TRY_AGAIN (WSATRY_AGAIN)
value TT_POLYGON_TYPE (24)
value TT_PRIM_CSPLINE (3)
value TT_PRIM_LINE (1)
value TT_PRIM_QSPLINE (2)
value TURKISH_CHARSET (162)
value TWOSTOPBITS (2)
value TXFS_RM_STATE_ACTIVE (2)
value TXFS_RM_STATE_NOT_STARTED (0)
value TXFS_RM_STATE_SHUTTING_DOWN (3)
value TXFS_RM_STATE_STARTING (1)
value UILANGUAGE_ENUMPROC (UILANGUAGE_ENUMPROCA)
value UIS_CLEAR (2)
value UIS_INITIALIZE (3)
value UIS_SET (1)
value UMS_VERSION (RTL_UMS_VERSION)
value UNLOAD_DLL_DEBUG_EVENT (7)
value UNLOCK_ELEMENT (1)
value UNWIND_CHAIN_LIMIT (32)
value UNWIND_HISTORY_TABLE_SIZE (12)
value UOI_FLAGS (1)
value UOI_HEAPSIZE (5)
value UOI_IO (6)
value UOI_NAME (2)
value UOI_TIMERPROC_EXCEPTION_SUPPRESSION (7)
value UOI_TYPE (3)
value UOI_USER_SID (4)
value URL_MK_LEGACY (0)
value URL_MK_NO_CANONICALIZE (2)
value URL_MK_UNIFORM (1)
value USER_DEFAULT_SCREEN_DPI (96)
value USER_MARSHAL_FC_BYTE (1)
value USER_MARSHAL_FC_CHAR (2)
value USER_MARSHAL_FC_DOUBLE (12)
value USER_MARSHAL_FC_FLOAT (10)
value USER_MARSHAL_FC_HYPER (11)
value USER_MARSHAL_FC_LONG (8)
value USER_MARSHAL_FC_SHORT (6)
value USER_MARSHAL_FC_SMALL (3)
value USER_MARSHAL_FC_ULONG (9)
value USER_MARSHAL_FC_USHORT (7)
value USER_MARSHAL_FC_USMALL (4)
value USER_MARSHAL_FC_WCHAR (5)
value VARCMP_EQ (1)
value VARCMP_GT (2)
value VARCMP_LT (0)
value VARCMP_NULL (3)
value VARIABLE_PITCH (2)
value VENDOR_ID_LENGTH (8)
value VERTRES (10)
value VERTSIZE (6)
value VER_AND (6)
value VER_CONDITION_MASK (7)
value VER_EQUAL (1)
value VER_GREATER (2)
value VER_GREATER_EQUAL (3)
value VER_LESS (4)
value VER_LESS_EQUAL (5)
value VER_NUM_BITS_PER_CONDITION_MASK (3)
value VER_OR (7)
value VIETNAMESE_CHARSET (163)
value VREFRESH (116)
value VS_FILE_INFO (RT_VERSION)
value VS_USER_DEFINED (100)
value VS_VERSION_INFO (1)
value VTA_BASELINE (TA_BASELINE)
value VTA_BOTTOM (TA_RIGHT)
value VTA_CENTER (TA_CENTER)
value VTA_LEFT (TA_BOTTOM)
value VTA_RIGHT (TA_TOP)
value VTA_TOP (TA_LEFT)
value VTDATEGRE_MAX (2958465)
value VT_HARDTYPE (VT_RESERVED)
value WAIT_IO_COMPLETION (STATUS_USER_APC)
value WAIT_TIMEOUT (258L)
value WARNING_IPSEC_MM_POLICY_PRUNED (13024L)
value WARNING_IPSEC_QM_POLICY_PRUNED (13025L)
value WAVERR_BASE (32)
value WAVE_FORMAT_PCM (1)
value WA_ACTIVE (1)
value WA_CLICKACTIVE (2)
value WA_INACTIVE (0)
value WB_ISDELIMITER (2)
value WB_LEFT (0)
value WB_RIGHT (1)
value WDK_NTDDI_VERSION (NTDDI_WIN10_NI)
value WGL_FONT_LINES (0)
value WGL_FONT_POLYGONS (1)
value WGL_SWAPMULTIPLE_MAX (16)
value WHEEL_DELTA (120)
value WHITEONBLACK (2)
value WHITE_BRUSH (0)
value WHITE_PEN (6)
value WH_CALLWNDPROC (4)
value WH_CALLWNDPROCRET (12)
value WH_CBT (5)
value WH_DEBUG (9)
value WH_FOREGROUNDIDLE (11)
value WH_GETMESSAGE (3)
value WH_JOURNALPLAYBACK (1)
value WH_JOURNALRECORD (0)
value WH_KEYBOARD (2)
value WH_KEYBOARD_LL (13)
value WH_MAX (14)
value WH_MAXHOOK (WH_MAX)
value WH_MINHOOK (WH_MIN)
value WH_MOUSE (7)
value WH_MOUSE_LL (14)
value WH_SHELL (10)
value WH_SYSMSGFILTER (6)
value WIM_CLOSE (MM_WIM_CLOSE)
value WIM_DATA (MM_WIM_DATA)
value WIM_OPEN (MM_WIM_OPEN)
value WIM_PROVIDER_HASH_SIZE (20)
value WINABLEAPI (DECLSPEC_IMPORT)
value WINADVAPI (DECLSPEC_IMPORT)
value WINAPI_FAMILY (WINAPI_FAMILY_DESKTOP_APP)
value WINAPI_FAMILY_APP (WINAPI_FAMILY_PC_APP)
value WINAPI_FAMILY_DESKTOP_APP (100)
value WINAPI_FAMILY_GAMES (6)
value WINAPI_FAMILY_PC_APP (2)
value WINAPI_FAMILY_PHONE_APP (3)
value WINAPI_FAMILY_SERVER (5)
value WINAPI_FAMILY_SYSTEM (4)
value WINAPI_INLINE (WINAPI)
value WINAPI_PARTITION_PHONE (WINAPI_PARTITION_PHONE_APP)
value WINBASEAPI (DECLSPEC_IMPORT)
value WINCOMMCTRLAPI (DECLSPEC_IMPORT)
value WINCOMMDLGAPI (DECLSPEC_IMPORT)
value WINDEVQUERYAPI (DECLSPEC_IMPORT)
value WINDING (2)
value WINGDIAPI (DECLSPEC_IMPORT)
value WININETINFO_OPTION_LOCK_HANDLE (65534)
value WINMMAPI (DECLSPEC_IMPORT)
value WINNORMALIZEAPI (DECLSPEC_IMPORT)
value WINPATHCCHAPI (WINBASEAPI)
value WINPERF_LOG_DEBUG (2)
value WINPERF_LOG_NONE (0)
value WINPERF_LOG_USER (1)
value WINPERF_LOG_VERBOSE (3)
value WINSHELLAPI (DECLSPEC_IMPORT)
value WINSOCK_API_LINKAGE (DECLSPEC_IMPORT)
value WINSPOOLAPI (DECLSPEC_IMPORT)
value WINSTORAGEAPI (DECLSPEC_IMPORT)
value WINSWDEVICEAPI (DECLSPEC_IMPORT)
value WINUSERAPI (DECLSPEC_IMPORT)
value WINVER (_WIN32_WINNT)
value WIZ_BODYCX (184)
value WIZ_BODYX (92)
value WIZ_CXBMP (80)
value WIZ_CXDLG (276)
value WIZ_CYDLG (140)
value WMSZ_BOTTOM (6)
value WMSZ_BOTTOMLEFT (7)
value WMSZ_BOTTOMRIGHT (8)
value WMSZ_LEFT (1)
value WMSZ_RIGHT (2)
value WMSZ_TOP (3)
value WMSZ_TOPLEFT (4)
value WMSZ_TOPRIGHT (5)
value WM_SETTINGCHANGE (WM_WININICHANGE)
value WNNC_NET_LANMAN (WNNC_NET_SMB)
value WN_ACCESS_DENIED (ERROR_ACCESS_DENIED)
value WN_ALREADY_CONNECTED (ERROR_ALREADY_ASSIGNED)
value WN_BAD_DEV_TYPE (ERROR_BAD_DEV_TYPE)
value WN_BAD_HANDLE (ERROR_INVALID_HANDLE)
value WN_BAD_LEVEL (ERROR_INVALID_LEVEL)
value WN_BAD_LOCALNAME (ERROR_BAD_DEVICE)
value WN_BAD_NETNAME (ERROR_BAD_NET_NAME)
value WN_BAD_PASSWORD (ERROR_INVALID_PASSWORD)
value WN_BAD_POINTER (ERROR_INVALID_ADDRESS)
value WN_BAD_PROFILE (ERROR_BAD_PROFILE)
value WN_BAD_PROVIDER (ERROR_BAD_PROVIDER)
value WN_BAD_USER (ERROR_BAD_USERNAME)
value WN_BAD_VALUE (ERROR_INVALID_PARAMETER)
value WN_CANCEL (ERROR_CANCELLED)
value WN_CANNOT_OPEN_PROFILE (ERROR_CANNOT_OPEN_PROFILE)
value WN_CONNECTED_OTHER_PASSWORD (ERROR_CONNECTED_OTHER_PASSWORD)
value WN_CONNECTED_OTHER_PASSWORD_DEFAULT (ERROR_CONNECTED_OTHER_PASSWORD_DEFAULT)
value WN_CONNECTION_CLOSED (ERROR_CONNECTION_UNAVAIL)
value WN_DEVICE_ALREADY_REMEMBERED (ERROR_DEVICE_ALREADY_REMEMBERED)
value WN_DEVICE_ERROR (ERROR_GEN_FAILURE)
value WN_DEVICE_IN_USE (ERROR_DEVICE_IN_USE)
value WN_EXTENDED_ERROR (ERROR_EXTENDED_ERROR)
value WN_FUNCTION_BUSY (ERROR_BUSY)
value WN_MORE_DATA (ERROR_MORE_DATA)
value WN_NET_ERROR (ERROR_UNEXP_NET_ERR)
value WN_NOT_AUTHENTICATED (ERROR_NOT_AUTHENTICATED)
value WN_NOT_CONNECTED (ERROR_NOT_CONNECTED)
value WN_NOT_CONTAINER (ERROR_NOT_CONTAINER)
value WN_NOT_INITIALIZING (ERROR_ALREADY_INITIALIZED)
value WN_NOT_LOGGED_ON (ERROR_NOT_LOGGED_ON)
value WN_NOT_SUPPORTED (ERROR_NOT_SUPPORTED)
value WN_NOT_VALIDATED (ERROR_NO_LOGON_SERVERS)
value WN_NO_ERROR (NO_ERROR)
value WN_NO_MORE_DEVICES (ERROR_NO_MORE_DEVICES)
value WN_NO_MORE_ENTRIES (ERROR_NO_MORE_ITEMS)
value WN_NO_NETWORK (ERROR_NO_NETWORK)
value WN_NO_NET_OR_BAD_PATH (ERROR_NO_NET_OR_BAD_PATH)
value WN_OPEN_FILES (ERROR_OPEN_FILES)
value WN_OUT_OF_MEMORY (ERROR_NOT_ENOUGH_MEMORY)
value WN_RETRY (ERROR_RETRY)
value WN_SUCCESS (NO_ERROR)
value WN_WINDOWS_ERROR (ERROR_UNEXP_NET_ERR)
value WOM_CLOSE (MM_WOM_CLOSE)
value WOM_DONE (MM_WOM_DONE)
value WOM_OPEN (MM_WOM_OPEN)
value WSABASEERR (10000)
value WSADESCRIPTION_LEN (256)
value WSAEACCES (10013L)
value WSAEADDRINUSE (10048L)
value WSAEADDRNOTAVAIL (10049L)
value WSAEAFNOSUPPORT (10047L)
value WSAEALREADY (10037L)
value WSAEBADF (10009L)
value WSAECANCELLED (10103L)
value WSAECONNABORTED (10053L)
value WSAECONNREFUSED (10061L)
value WSAECONNRESET (10054L)
value WSAEDESTADDRREQ (10039L)
value WSAEDISCON (10101L)
value WSAEDQUOT (10069L)
value WSAEFAULT (10014L)
value WSAEHOSTDOWN (10064L)
value WSAEHOSTUNREACH (10065L)
value WSAEINPROGRESS (10036L)
value WSAEINTR (10004L)
value WSAEINVAL (10022L)
value WSAEINVALIDPROCTABLE (10104L)
value WSAEINVALIDPROVIDER (10105L)
value WSAEISCONN (10056L)
value WSAELOOP (10062L)
value WSAEMFILE (10024L)
value WSAEMSGSIZE (10040L)
value WSAENAMETOOLONG (10063L)
value WSAENETDOWN (10050L)
value WSAENETRESET (10052L)
value WSAENETUNREACH (10051L)
value WSAENOBUFS (10055L)
value WSAENOMORE (10102L)
value WSAENOPROTOOPT (10042L)
value WSAENOTCONN (10057L)
value WSAENOTEMPTY (10066L)
value WSAENOTSOCK (10038L)
value WSAEOPNOTSUPP (10045L)
value WSAEPFNOSUPPORT (10046L)
value WSAEPROCLIM (10067L)
value WSAEPROTONOSUPPORT (10043L)
value WSAEPROTOTYPE (10041L)
value WSAEPROVIDERFAILEDINIT (10106L)
value WSAEREFUSED (10112L)
value WSAEREMOTE (10071L)
value WSAESHUTDOWN (10058L)
value WSAESOCKTNOSUPPORT (10044L)
value WSAESTALE (10070L)
value WSAETIMEDOUT (10060L)
value WSAETOOMANYREFS (10059L)
value WSAEUSERS (10068L)
value WSAEVENT (HANDLE)
value WSAEWOULDBLOCK (10035L)
value WSAHOST_NOT_FOUND (11001L)
value WSANOTINITIALISED (10093L)
value WSANO_ADDRESS (WSANO_DATA)
value WSANO_DATA (11004L)
value WSANO_RECOVERY (11003L)
value WSAOVERLAPPED (OVERLAPPED)
value WSAPROTOCOL_LEN (255)
value WSASERVICE_NOT_FOUND (10108L)
value WSASYSCALLFAILURE (10107L)
value WSASYSNOTREADY (10091L)
value WSASYS_STATUS_LEN (128)
value WSATRY_AGAIN (11002L)
value WSATYPE_NOT_FOUND (10109L)
value WSAVERNOTSUPPORTED (10092L)
value WSA_E_CANCELLED (10111L)
value WSA_E_NO_MORE (10110L)
value WSA_IPSEC_NAME_POLICY_ERROR (11033L)
value WSA_QOS_ADMISSION_FAILURE (11010L)
value WSA_QOS_BAD_OBJECT (11013L)
value WSA_QOS_BAD_STYLE (11012L)
value WSA_QOS_EFILTERCOUNT (11021L)
value WSA_QOS_EFILTERSTYLE (11019L)
value WSA_QOS_EFILTERTYPE (11020L)
value WSA_QOS_EFLOWCOUNT (11023L)
value WSA_QOS_EFLOWDESC (11026L)
value WSA_QOS_EFLOWSPEC (11017L)
value WSA_QOS_EOBJLENGTH (11022L)
value WSA_QOS_EPOLICYOBJ (11025L)
value WSA_QOS_EPROVSPECBUF (11018L)
value WSA_QOS_EPSFILTERSPEC (11028L)
value WSA_QOS_EPSFLOWSPEC (11027L)
value WSA_QOS_ESDMODEOBJ (11029L)
value WSA_QOS_ESERVICETYPE (11016L)
value WSA_QOS_ESHAPERATEOBJ (11030L)
value WSA_QOS_EUNKOWNPSOBJ (11024L)
value WSA_QOS_GENERIC_ERROR (11015L)
value WSA_QOS_NO_RECEIVERS (11008L)
value WSA_QOS_NO_SENDERS (11007L)
value WSA_QOS_POLICY_FAILURE (11011L)
value WSA_QOS_RECEIVERS (11005L)
value WSA_QOS_REQUEST_CONFIRMED (11009L)
value WSA_QOS_RESERVED_PETYPE (11031L)
value WSA_QOS_SENDERS (11006L)
value WSA_QOS_TRAFFIC_CTRL_ERROR (11014L)
value WSA_SECURE_HOST_NOT_FOUND (11032L)
value WS_ICONIC (WS_MINIMIZE)
value WS_SIZEBOX (WS_THICKFRAME)
value WS_TILED (WS_OVERLAPPED)
value WS_TILEDWINDOW (WS_OVERLAPPEDWINDOW)
value XST_ADVACKRCVD (13)
value XST_ADVDATAACKRCVD (16)
value XST_ADVDATASENT (15)
value XST_ADVSENT (11)
value XST_CONNECTED (2)
value XST_DATARCVD (6)
value XST_EXECACKRCVD (10)
value XST_EXECSENT (9)
value XST_INCOMPLETE (1)
value XST_NULL (0)
value XST_POKEACKRCVD (8)
value XST_POKESENT (7)
value XST_REQSENT (5)
value XST_UNADVACKRCVD (14)
value XST_UNADVSENT (12)
value XTYP_SHIFT (4)
value ZAWPROXYAPI (DECLSPEC_IMPORT)
value ZERO_PADDING (3)
value _ACRTIMP_ALT (_ACRTIMP)
value _ARGMAX (100)
value _ARM_WINAPI_PARTITION_DESKTOP_SDK_AVAILABLE (1)
value _ASSEMBLY_DLL_REDIRECTION_DETAILED_INFORMATION (_ASSEMBLY_FILE_DETAILED_INFORMATION)
value _CRT_BUILD_DESKTOP_APP (1)
value _CRT_FUNCTIONS_REQUIRED (1)
value _CRT_INTERNAL_NONSTDC_NAMES (1)
value _CRT_INT_MAX (2147483647)
value _CRT_PACKING (8)
value _CRT_SECURE_CPP_OVERLOAD_SECURE_NAMES (1)
value _CRT_SECURE_CPP_OVERLOAD_SECURE_NAMES_MEMORY (0)
value _CRT_SECURE_CPP_OVERLOAD_STANDARD_NAMES (0)
value _CRT_SECURE_CPP_OVERLOAD_STANDARD_NAMES_COUNT (0)
value _CRT_SECURE_CPP_OVERLOAD_STANDARD_NAMES_MEMORY (0)
value _CRT_USE_CONFORMING_ANNEX_K_TIME (0)
value _HAS_EXCEPTIONS (1)
value _HAS_NODISCARD (0)
value _INTEGRAL_MAX_BITS (64)
value _IOB_ENTRIES (3)
value _MAX_DIR (256)
value _MAX_DRIVE (3)
value _MAX_ENV (32767)
value _MAX_EXT (256)
value _MAX_FNAME (256)
value _MAX_PATH (260)
value _MM_HINT_NTA (0)
value _MSC_BUILD (1)
value _MSC_EXTENSIONS (1)
value _MSC_FULL_VER (192000000)
value _MSC_VER (1920)
value _MSVC_EXECUTION_CHARACTER_SET (65001)
value _NFILE (_NSTREAM_)
value _NLSCMPERROR (_CRT_INT_MAX)
value _NSTREAM_ (512)
value _OUT_TO_DEFAULT (0)
value _OUT_TO_MSGBOX (2)
value _OUT_TO_STDERR (1)
value _O_RAW (_O_BINARY)
value _REPORT_ERRMODE (3)
value _RPC_HTTP_TRANSPORT_CREDENTIALS (_RPC_HTTP_TRANSPORT_CREDENTIALS_A)
value _SAL_VERSION (20)
value _SEC_WINNT_AUTH_IDENTITY (_SEC_WINNT_AUTH_IDENTITY_A)
value _SS_MAXSIZE (128)
value _STRALIGN_USE_SECURE_CRT (1)
value _SYS_OPEN (20)
value _TMP_MAX_S (TMP_MAX)
value _USE_ATTRIBUTES_FOR_SAL (0)
value _USE_DECLSPECS_FOR_SAL (0)
value _VCRT_COMPILER_PREPROCESSOR (1)
value __ATOMIC_ACQUIRE (2)
value __ATOMIC_ACQ_REL (4)
value __ATOMIC_CONSUME (1)
value __ATOMIC_RELAXED (0)
value __ATOMIC_RELEASE (3)
value __ATOMIC_SEQ_CST (5)
value __BIGGEST_ALIGNMENT__ (16)
value __BITINT_MAXWIDTH__ (128)
value __BOOL_WIDTH__ (8)
value __BYTE_ORDER__ (__ORDER_LITTLE_ENDIAN__)
value __CHAR_BIT__ (8)
value __CLANG_ATOMIC_BOOL_LOCK_FREE (2)
value __CLANG_ATOMIC_CHAR_LOCK_FREE (2)
value __CLANG_ATOMIC_INT_LOCK_FREE (2)
value __CLANG_ATOMIC_LLONG_LOCK_FREE (2)
value __CLANG_ATOMIC_LONG_LOCK_FREE (2)
value __CLANG_ATOMIC_POINTER_LOCK_FREE (2)
value __CLANG_ATOMIC_SHORT_LOCK_FREE (2)
value __CLANG_ATOMIC_WCHAR_T_LOCK_FREE (2)
value __CONSTANT_CFSTRINGS__ (1)
value __CRTDECL (__CLRCALL_PURE_OR_CDECL)
value __DBL_DECIMAL_DIG__ (17)
value __DBL_DIG__ (15)
value __DBL_HAS_DENORM__ (1)
value __DBL_HAS_INFINITY__ (1)
value __DBL_HAS_QUIET_NAN__ (1)
value __DBL_MANT_DIG__ (53)
value __DBL_MAX_EXP__ (1024)
value __DECIMAL_DIG__ (__LDBL_DECIMAL_DIG__)
value __FINITE_MATH_ONLY__ (0)
value __FLT_DECIMAL_DIG__ (9)
value __FLT_DIG__ (6)
value __FLT_HAS_DENORM__ (1)
value __FLT_HAS_INFINITY__ (1)
value __FLT_HAS_QUIET_NAN__ (1)
value __FLT_MANT_DIG__ (24)
value __FLT_MAX_EXP__ (128)
value __FLT_RADIX__ (2)
value __FXSR__ (1)
value __GCC_ASM_FLAG_OUTPUTS__ (1)
value __GOT_SECURE_LIB__ (__STDC_SECURE_LIB__)
value __INTMAX_C_SUFFIX__ (LL)
value __INTMAX_MAX__ (9223372036854775807LL)
value __INTMAX_WIDTH__ (64)
value __INTPTR_MAX__ (9223372036854775807LL)
value __INTPTR_WIDTH__ (64)
value __INT_MAX__ (2147483647)
value __INT_WIDTH__ (32)
value __LDBL_DECIMAL_DIG__ (17)
value __LDBL_DIG__ (15)
value __LDBL_HAS_DENORM__ (1)
value __LDBL_HAS_INFINITY__ (1)
value __LDBL_HAS_QUIET_NAN__ (1)
value __LDBL_MANT_DIG__ (53)
value __LDBL_MAX_EXP__ (1024)
value __LITTLE_ENDIAN__ (1)
value __LLONG_WIDTH__ (64)
value __LONG_LONG_MAX__ (9223372036854775807LL)
value __LONG_MAX__ (2147483647L)
value __LONG_WIDTH__ (32)
value __MMX__ (1)
value __NO_INLINE__ (1)
value __NO_MATH_INLINES (1)
value __OBJC_BOOL_IS_BOOL (0)
value __OPENCL_MEMORY_SCOPE_ALL_SVM_DEVICES (3)
value __OPENCL_MEMORY_SCOPE_DEVICE (2)
value __OPENCL_MEMORY_SCOPE_SUB_GROUP (4)
value __OPENCL_MEMORY_SCOPE_WORK_GROUP (1)
value __OPENCL_MEMORY_SCOPE_WORK_ITEM (0)
value __ORDER_BIG_ENDIAN__ (4321)
value __ORDER_LITTLE_ENDIAN__ (1234)
value __ORDER_PDP_ENDIAN__ (3412)
value __PIC__ (2)
value __POINTER_WIDTH__ (64)
value __PRAGMA_REDEFINE_EXTNAME (1)
value __PTRDIFF_MAX__ (9223372036854775807LL)
value __PTRDIFF_WIDTH__ (64)
value __REQUIRED_RPCNDR_H_VERSION__ (501)
value __REQUIRED_RPCSAL_H_VERSION__ (100)
value __SAL_H_FULL_VER (140050727)
value __SAL_H_VERSION (180000000)
value __SCHAR_MAX__ (127)
value __SEG_FS (1)
value __SEG_GS (1)
value __SHRT_MAX__ (32767)
value __SHRT_WIDTH__ (16)
value __SIG_ATOMIC_MAX__ (2147483647)
value __SIG_ATOMIC_WIDTH__ (32)
value __SIZEOF_DOUBLE__ (8)
value __SIZEOF_FLOAT__ (4)
value __SIZEOF_INT__ (4)
value __SIZEOF_LONG_DOUBLE__ (8)
value __SIZEOF_LONG_LONG__ (8)
value __SIZEOF_LONG__ (4)
value __SIZEOF_POINTER__ (8)
value __SIZEOF_PTRDIFF_T__ (8)
value __SIZEOF_SHORT__ (2)
value __SIZEOF_SIZE_T__ (8)
value __SIZEOF_WCHAR_T__ (2)
value __SIZEOF_WINT_T__ (2)
value __SIZE_MAX__ (18446744073709551615ULL)
value __SIZE_WIDTH__ (64)
value __SPECSTRINGS_STRICT_LEVEL (1)
value __SSE_MATH__ (1)
value __SSE__ (1)
value __STDC_HOSTED__ (1)
value __STDC_NO_THREADS__ (1)
value __STDC_SECURE_LIB__ (200411L)
value __STDC_VERSION__ (201710L)
value __STDC_WANT_SECURE_LIB__ (1)
value __UINTMAX_C_SUFFIX__ (ULL)
value __UINTMAX_MAX__ (18446744073709551615ULL)
value __UINTMAX_WIDTH__ (64)
value __UINTPTR_MAX__ (18446744073709551615ULL)
value __UINTPTR_WIDTH__ (64)
value __WCHAR_MAX__ (65535)
value __WCHAR_UNSIGNED__ (1)
value __WCHAR_WIDTH__ (16)
value __WINT_MAX__ (65535)
value __WINT_UNSIGNED__ (1)
value __WINT_WIDTH__ (16)

