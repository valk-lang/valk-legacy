

fn write(fd: i32, data: ptr, length: uint);
