
fn malloc(size: uint) ptr;
fn write(fd: i32, data: ptr, length: uint);
