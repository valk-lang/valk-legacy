
value INFINITE (4294967295)
value EAGAIN (536870918)
value EWOULDBLOCK (536871039)
value SOCK_STREAM (1)

value SOL_SOCKET (65535)
value SO_REUSEADDR (4)
value SO_RCVTIMEO (4102)

value AF_INET (2)
value AF_UNIX (1)

value AI_PASSIVE (1)
value AI_CANONNAME (2)
value AI_NUMERICHOST (4)

value POLLIN (768)
value POLLOUT (16)
value POLLERR (1)
value POLLHUP (2)

// WSA
value WSAEWOULDBLOCK (10035)
value WSAENOBUFS (10055)
value FIONBIO (2148034174)

value O_RDONLY (0)
value O_WRONLY (1)
value O_RDWR (2)

value O_APPEND (8)
value O_CREATE (256)
value O_TRUNC (512)
value O_EXCL (1024)
value O_SYNC (4096)

value S_IFDIR (16384)
value S_IFREG (32768)
value S_IFMT (126976)

value INVALID_FILE_ATTRIBUTES (4294967295)
value FILE_ATTRIBUTE_ARCHIVE (32)
value FILE_ATTRIBUTE_DIRECTORY (16)
value FILE_ATTRIBUTE_HIDDEN (2)
value FILE_ATTRIBUTE_NORMAL (128)
value FILE_ATTRIBUTE_READONLY (1)
value FILE_ATTRIBUTE_SYSTEM (4)
