
value EINTR (4)
value EAGAIN (11)
value EWOULDBLOCK (11)
value EINVAL (22)

value SOCK_STREAM (1)
value SOCK_NONBLOCK (2048)

value SOL_SOCKET (1)
value SOL_TCP (6)
value SO_REUSEADDR (2)
value SO_RCVTIMEO (20)

value AF_INET (2)
value AF_UNIX (1)

value AI_PASSIVE (1)
value AI_CANONNAME (2)
value AI_NUMERICHOST (4)

value POLLIN (1)
value POLLOUT (4)
value POLLERR (8)
value POLLHUP (16)
value POLLRDHUP (8192)

value EPOLLERR (8)
value EPOLLET (-2147483648)
value EPOLLHUP (16)
value EPOLLIN (1)
value EPOLLMSG (1024)
value EPOLLONESHOT (1073741824)
value EPOLLOUT (4)
value EPOLLPRI (2)
value EPOLLRDBAND (128)
value EPOLLRDHUP (8192)
value EPOLLRDNORM (64)
value EPOLLWRBAND (512)
value EPOLLWRNORM (256)
value EPOLL_CLOEXEC (524288)
value EPOLL_CTL_ADD (1)
value EPOLL_CTL_DEL (2)
value EPOLL_CTL_MOD (3)
value EPOLL_NONBLOCK (2048)

value O_RDONLY (0)
value O_RDWR (2)
value O_WRONLY (1)
//
value O_CREATE (64)
value O_EXCL (128)
value O_TRUNC (512)
value O_APPEND (1024)
value O_NONBLOCK (2048)
value O_SYNC (1052672)

value S_IFDIR (16384)
value S_IFREG (32768)
value S_IFMT (61440)