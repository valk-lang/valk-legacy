
value EAGAIN (35)
value SOCK_STREAM (1)
value F_GETFL (3)
value F_SETFL (4)
value O_NONBLOCK (4)

value SOL_SOCKET (65535)
value SO_REUSEADDR (4)
value SO_RCVTIMEO (4102)

value AF_INET (2)
value AF_UNIX (1)

value AI_PASSIVE (1)
value AI_CANONNAME (2)
value AI_NUMERICHOST (4)

value POLLIN (1)
value POLLOUT (4)
value POLLERR (8)
value POLLHUP (16)
value POLLRDHUP (8192)

value O_RDONLY (0)
value O_RDWR (2)
value O_WRONLY (1)

value O_APPEND (8)
value O_CREATE (512)
value O_EXCL (2048)
value O_SYNC (128)
value O_TRUNC (1024)

value S_IFDIR (16384)
value S_IFREG (32768)
value S_IFMT (61440)
