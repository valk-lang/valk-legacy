
struct libc_jmp_buf {
    data: inline [ptr, 5]
}

struct libc_stat {
    st_dev: uint
    st_ino: uint
    st_nlink: uint
    st_mode: u32
    st_uid: u32
    st_gid: u32
    __pad0: u32
    st_rdev: uint
    st_size: int
    st_blksize: int
    st_blocks: int // Number 512-byte blocks allocated
    st_atime: uint
    st_atime_nsec: uint
    st_mtime: uint
    st_mtime_nsec: uint
    st_ctime: uint
    st_ctime_nsec: uint
    __unused_1: int
    __unused_2: int
    __unused_3: int
}

struct libc_timespec {
    tv_sec: int // seconds
    tv_nsec: int // nanoseconds
}

struct libc_timeval {
    tv_sec: int // seconds
    tv_usec: int // microseconds
}

struct libc_pollfd {
    fd: int // SOCKET (aka. HANDLE)
    events: i16  // detect events
    revents: i16 // detected events
}

struct libc_addrinfo {
    ai_flags: i32
    ai_family: i32
    ai_socktype: i32
    ai_protocol: i32
    ai_addrlen: uint
    ai_canonname: cstring
    ai_addr: libc_sockaddr
    ai_next: ?libc_addrinfo
}

struct libc_sockaddr {
    sa_family: u16
    sa_data_1: u32
    sa_data_2: u32
    sa_data_3: u32
    sa_data_4: u16
}

//struct libc_sockaddr_in {
//    sin_family: i16
//    sin_port: u16
//    sin_addr: .libc_in_addr
//    sin_zero: .u8[8]
//}

struct libc_in_addr {
    S_addr: u32
}

//struct WSADATA {
//    wVersion: u16
//    wHighVersion: u16
//
//    // 64-bit fields
//    iMaxSockets: u16
//    iMaxUdpDg: u16
//    lpVendorInfo: cstring
//    szDescription: inline u8[257] // WSADESCRIPTION_LEN + 1
//    szSystemStatus: inline u8[257]
//
//    // 32-bit fields
//    //szDescription: inline u8[257]
//    //szSystemStatus: inline u8[257]
//    //iMaxSockets: u16
//    //iMaxUdpDg: u16
//    //lpVendorInfo: cstring
//}

struct libc_timezone {
    tz_minuteswest: i32 // Minutes west of GMT
    tz_dsttime: i32 // Nonzero if DST is ever in effect
}

struct WIN32_FIND_DATAA {
    dwFileAttributes: i32
    ftCreationTime: inline FILETIME
    ftLastAccessTime: inline FILETIME
    ftLastWriteTime: inline FILETIME
    nFileSizeHigh: i32
    nFileSizeLow: i32
    dwReserved0: i32
    dwReserved1: i32
    cFileName: inline [i8, 260]
    cAlternateFileName: inline [i8, 14]
    dwFileType: i32 // Obsolete. Do not use.
    dwCreatorType: i32 // Obsolete. Do not use
    wFinderFlags: i16 // Obsolete. Do not use
}

struct FILETIME {
    dwLowDateTime: i32
    dwHighDateTime: i32
}

struct WSPUPCALLTABLE {
    lpWPUCloseEvent: ptr
    lpWPUCloseSocketHandle: ptr
    lpWPUCreateEvent: ptr
    lpWPUCreateSocketHandle: ptr
    lpWPUFDIsSet: ptr
    lpWPUGetProviderPath: ptr
    lpWPUModifyIFSHandle: ptr
    lpWPUPostMessage: ptr
    lpWPUQueryBlockingCallback: ptr
    lpWPUQuerySocketHandleContext: ptr
    lpWPUQueueApc: ptr
    lpWPUResetEvent: ptr
    lpWPUSetEvent: ptr
    lpWPUOpenCurrentThread: ptr
    lpWPUCloseThread: ptr
}

struct WSPPROC_TABLE {
    lpWSPAccept: ptr
    lpWSPAddressToString: ptr
    lpWSPAsyncSelect: ptr
    lpWSPBind: ptr
    lpWSPCancelBlockingCall: ptr
    lpWSPCleanup: ptr
    lpWSPCloseSocket: ptr
    lpWSPConnect: ptr
    lpWSPDuplicateSocket: ptr
    lpWSPEnumNetworkEvents: ptr
    lpWSPEventSelect: ptr
    lpWSPGetOverlappedResult: ptr
    lpWSPGetPeerName: ptr
    lpWSPGetSockName: ptr
    lpWSPGetSockOpt: ptr
    lpWSPGetQOSByName: ptr
    lpWSPIoctl: ptr
    lpWSPJoinLeaf: ptr
    lpWSPListen: ptr
    lpWSPRecv: ptr
    lpWSPRecvDisconnect: ptr
    lpWSPRecvFrom: ptr
    lpWSPSelect: ptr
    lpWSPSend: ptr
    lpWSPSendDisconnect: ptr
    lpWSPSendTo: ptr
    lpWSPSetSockOpt: ptr
    lpWSPShutdown: ptr
    lpWSPSocket: ptr
    lpWSPStringToAddress: ptr
}

struct _GUID {
  Data1: u32
  Data2: u16
  Data3: u16
  Data4: u64 // or .u8[8]
}

// struct WSAPROTOCOLCHAIN {
//   ChainLen: i32
//   ChainEntries: .u32[7] //DWORD ChainEntries[MAX_PROTOCOL_CHAIN]
// }

// struct WSAPROTOCOL_INFOA {
//   dwServiceFlags1: u32
//   dwServiceFlags2: u32
//   dwServiceFlags3: u32
//   dwServiceFlags4: u32
//   dwProviderFlags: u32
//   ProviderId: ._GUID
//   dwCatalogEntryId: u32
//   ProtocolChain: .WSAPROTOCOLCHAIN
//   iVersion: i32
//   iAddressFamily: i32
//   iMaxSockAddr: i32
//   iMinSockAddr: i32
//   iSocketType: i32
//   iProtocol: i32
//   iProtocolMaxOffset: i32
//   iNetworkByteOrder: i32
//   iSecurityScheme: i32
//   dwMessageSize: u32
//   dwProviderReserved: u32
//   szProtocol: .u8[256] //CHAR szProtocol[WSAPROTOCOL_LEN + 1]
// }

// struct WSPDATA {
//   wVersion: u16
//   wHighVersion: u16
//   szDescription: .u16[256] //WCHAR szDescription[WSPDESCRIPTION_LEN + 1]
// }
