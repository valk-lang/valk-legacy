
value AF_ALG (PF_ALG)
value AF_APPLETALK (PF_APPLETALK)
value AF_ASH (PF_ASH)
value AF_ATMPVC (PF_ATMPVC)
value AF_ATMSVC (PF_ATMSVC)
value AF_BLUETOOTH (PF_BLUETOOTH)
value AF_BRIDGE (PF_BRIDGE)
value AF_CAIF (PF_CAIF)
value AF_CAN (PF_CAN)
value AF_ECONET (PF_ECONET)
value AF_FILE (PF_FILE)
value AF_IB (PF_IB)
value AF_INET (PF_INET)
value AF_IPX (PF_IPX)
value AF_IRDA (PF_IRDA)
value AF_ISDN (PF_ISDN)
value AF_IUCV (PF_IUCV)
value AF_KCM (PF_KCM)
value AF_KEY (PF_KEY)
value AF_LLC (PF_LLC)
value AF_LOCAL (PF_LOCAL)
value AF_MAX (PF_MAX)
value AF_MCTP (PF_MCTP)
value AF_MPLS (PF_MPLS)
value AF_NETBEUI (PF_NETBEUI)
value AF_NETLINK (PF_NETLINK)
value AF_NETROM (PF_NETROM)
value AF_NFC (PF_NFC)
value AF_PACKET (PF_PACKET)
value AF_PHONET (PF_PHONET)
value AF_PPPOX (PF_PPPOX)
value AF_QIPCRTR (PF_QIPCRTR)
value AF_RDS (PF_RDS)
value AF_ROSE (PF_ROSE)
value AF_ROUTE (PF_ROUTE)
value AF_RXRPC (PF_RXRPC)
value AF_SECURITY (PF_SECURITY)
value AF_SMC (PF_SMC)
value AF_SNA (PF_SNA)
value AF_TIPC (PF_TIPC)
value AF_UNIX (PF_UNIX)
value AF_UNSPEC (PF_UNSPEC)
value AF_VSOCK (PF_VSOCK)
value AF_WANPIPE (PF_WANPIPE)
value AF_XDP (PF_XDP)
value AIO_PRIO_DELTA_MAX (20)
value BIG_ENDIAN (__BIG_ENDIAN)
value BUFSIZ (8192)
value BYTE_ORDER (__BYTE_ORDER)
value DELAYTIMER_MAX (2147483647)
value DT_BLK (DT_BLK)
value DT_CHR (DT_CHR)
value DT_DIR (DT_DIR)
value DT_FIFO (DT_FIFO)
value DT_LNK (DT_LNK)
value DT_REG (DT_REG)
value DT_SOCK (DT_SOCK)
value DT_UNKNOWN (DT_UNKNOWN)
value DT_WHT (DT_WHT)
value EACCES (13)
value EADDRINUSE (98)
value EADDRNOTAVAIL (99)
value EADV (68)
value EAFNOSUPPORT (97)
value EAGAIN (11)
value EALREADY (114)
value EBADE (52)
value EBADF (9)
value EBADFD (77)
value EBADMSG (74)
value EBADR (53)
value EBADRQC (56)
value EBADSLT (57)
value EBFONT (59)
value EBUSY (16)
value ECANCELED (125)
value ECHILD (10)
value ECHRNG (44)
value ECOMM (70)
value ECONNABORTED (103)
value ECONNREFUSED (111)
value ECONNRESET (104)
value EDEADLK (35)
value EDEADLOCK (EDEADLK)
value EDESTADDRREQ (89)
value EDOM (33)
value EDOTDOT (73)
value EDQUOT (122)
value EEXIST (17)
value EFAULT (14)
value EFBIG (27)
value EHOSTDOWN (112)
value EHOSTUNREACH (113)
value EHWPOISON (133)
value EIDRM (43)
value EILSEQ (84)
value EINPROGRESS (115)
value EINTR (4)
value EINVAL (22)
value EIO (5)
value EISCONN (106)
value EISDIR (21)
value EISNAM (120)
value EKEYEXPIRED (127)
value EKEYREJECTED (129)
value EKEYREVOKED (128)
value ELIBACC (79)
value ELIBBAD (80)
value ELIBEXEC (83)
value ELIBMAX (82)
value ELIBSCN (81)
value ELNRNG (48)
value ELOOP (40)
value EMEDIUMTYPE (124)
value EMFILE (24)
value EMLINK (31)
value EMSGSIZE (90)
value EMULTIHOP (72)
value ENAMETOOLONG (36)
value ENAVAIL (119)
value ENETDOWN (100)
value ENETRESET (102)
value ENETUNREACH (101)
value ENFILE (23)
value ENOANO (55)
value ENOBUFS (105)
value ENOCSI (50)
value ENODATA (61)
value ENODEV (19)
value ENOENT (2)
value ENOEXEC (8)
value ENOKEY (126)
value ENOLCK (37)
value ENOLINK (67)
value ENOMEDIUM (123)
value ENOMEM (12)
value ENOMSG (42)
value ENONET (64)
value ENOPKG (65)
value ENOPROTOOPT (92)
value ENOSPC (28)
value ENOSR (63)
value ENOSTR (60)
value ENOSYS (38)
value ENOTBLK (15)
value ENOTCONN (107)
value ENOTDIR (20)
value ENOTEMPTY (39)
value ENOTNAM (118)
value ENOTRECOVERABLE (131)
value ENOTSOCK (88)
value ENOTSUP (EOPNOTSUPP)
value ENOTTY (25)
value ENOTUNIQ (76)
value ENXIO (6)
value EOPNOTSUPP (95)
value EOVERFLOW (75)
value EOWNERDEAD (130)
value EPERM (1)
value EPFNOSUPPORT (96)
value EPIPE (32)
value EPOLLERR (EPOLLERR)
value EPOLLET (EPOLLET)
value EPOLLEXCLUSIVE (EPOLLEXCLUSIVE)
value EPOLLHUP (EPOLLHUP)
value EPOLLIN (EPOLLIN)
value EPOLLMSG (EPOLLMSG)
value EPOLLONESHOT (EPOLLONESHOT)
value EPOLLOUT (EPOLLOUT)
value EPOLLPRI (EPOLLPRI)
value EPOLLRDBAND (EPOLLRDBAND)
value EPOLLRDHUP (EPOLLRDHUP)
value EPOLLRDNORM (EPOLLRDNORM)
value EPOLLWAKEUP (EPOLLWAKEUP)
value EPOLLWRBAND (EPOLLWRBAND)
value EPOLLWRNORM (EPOLLWRNORM)
value EPOLL_CLOEXEC (EPOLL_CLOEXEC)
value EPOLL_CTL_ADD (1)
value EPOLL_CTL_DEL (2)
value EPOLL_CTL_MOD (3)
value EPROTO (71)
value EPROTONOSUPPORT (93)
value EPROTOTYPE (91)
value ERANGE (34)
value EREMCHG (78)
value EREMOTE (66)
value EREMOTEIO (121)
value ERESTART (85)
value ERFKILL (132)
value EROFS (30)
value ESHUTDOWN (108)
value ESOCKTNOSUPPORT (94)
value ESPIPE (29)
value ESRCH (3)
value ESRMNT (69)
value ESTALE (116)
value ESTRPIPE (86)
value ETIME (62)
value ETIMEDOUT (110)
value ETOOMANYREFS (109)
value ETXTBSY (26)
value EUCLEAN (117)
value EUNATCH (49)
value EUSERS (87)
value EWOULDBLOCK (EAGAIN)
value EXDEV (18)
value EXFULL (54)
value FAPPEND (O_APPEND)
value FASYNC (O_ASYNC)
value FD_CLOEXEC (1)
value FD_SETSIZE (__FD_SETSIZE)
value FFSYNC (O_FSYNC)
value FILENAME_MAX (4096)
value FNDELAY (O_NDELAY)
value FNONBLOCK (O_NONBLOCK)
value FOPEN_MAX (16)
value F_DUPFD (0)
value F_DUPFD_CLOEXEC (1030)
value F_EXLCK (4)
value F_GETFD (1)
value F_GETFL (3)
value F_GETLK (5)
value F_GETOWN (__F_GETOWN)
value F_LOCK (1)
value F_OK (0)
value F_RDLCK (0)
value F_SETFD (2)
value F_SETFL (4)
value F_SETLK (6)
value F_SETLKW (7)
value F_SETOWN (__F_SETOWN)
value F_SHLCK (8)
value F_TEST (3)
value F_TLOCK (2)
value F_ULOCK (0)
value F_UNLCK (2)
value F_WRLCK (1)
value HOST_NAME_MAX (64)
value HOST_NOT_FOUND (1)
value INET_ADDRSTRLEN (16)
value IN_CLASSA_MAX (128)
value IN_CLASSA_NSHIFT (24)
value IN_CLASSB_MAX (65536)
value IN_CLASSB_NSHIFT (16)
value IN_CLASSC_NSHIFT (8)
value IN_LOOPBACKNET (127)
value IPPORT_RESERVED (1024)
value IPPROTO_AH (IPPROTO_AH)
value IPPROTO_BEETPH (IPPROTO_BEETPH)
value IPPROTO_COMP (IPPROTO_COMP)
value IPPROTO_DCCP (IPPROTO_DCCP)
value IPPROTO_DSTOPTS (IPPROTO_DSTOPTS)
value IPPROTO_EGP (IPPROTO_EGP)
value IPPROTO_ENCAP (IPPROTO_ENCAP)
value IPPROTO_ESP (IPPROTO_ESP)
value IPPROTO_ETHERNET (IPPROTO_ETHERNET)
value IPPROTO_FRAGMENT (IPPROTO_FRAGMENT)
value IPPROTO_GRE (IPPROTO_GRE)
value IPPROTO_HOPOPTS (IPPROTO_HOPOPTS)
value IPPROTO_ICMP (IPPROTO_ICMP)
value IPPROTO_IDP (IPPROTO_IDP)
value IPPROTO_IGMP (IPPROTO_IGMP)
value IPPROTO_IP (IPPROTO_IP)
value IPPROTO_IPIP (IPPROTO_IPIP)
value IPPROTO_MH (IPPROTO_MH)
value IPPROTO_MPLS (IPPROTO_MPLS)
value IPPROTO_MPTCP (IPPROTO_MPTCP)
value IPPROTO_MTP (IPPROTO_MTP)
value IPPROTO_NONE (IPPROTO_NONE)
value IPPROTO_PIM (IPPROTO_PIM)
value IPPROTO_PUP (IPPROTO_PUP)
value IPPROTO_RAW (IPPROTO_RAW)
value IPPROTO_ROUTING (IPPROTO_ROUTING)
value IPPROTO_RSVP (IPPROTO_RSVP)
value IPPROTO_SCTP (IPPROTO_SCTP)
value IPPROTO_TCP (IPPROTO_TCP)
value IPPROTO_TP (IPPROTO_TP)
value IPPROTO_UDP (IPPROTO_UDP)
value IPPROTO_UDPLITE (IPPROTO_UDPLITE)
value IP_ADD_MEMBERSHIP (35)
value IP_ADD_SOURCE_MEMBERSHIP (39)
value IP_BIND_ADDRESS_NO_PORT (24)
value IP_BLOCK_SOURCE (38)
value IP_CHECKSUM (23)
value IP_DEFAULT_MULTICAST_LOOP (1)
value IP_DEFAULT_MULTICAST_TTL (1)
value IP_DROP_MEMBERSHIP (36)
value IP_DROP_SOURCE_MEMBERSHIP (40)
value IP_FREEBIND (15)
value IP_HDRINCL (3)
value IP_IPSEC_POLICY (16)
value IP_MAX_MEMBERSHIPS (20)
value IP_MINTTL (21)
value IP_MSFILTER (41)
value IP_MTU (14)
value IP_MTU_DISCOVER (10)
value IP_MULTICAST_ALL (49)
value IP_MULTICAST_IF (32)
value IP_MULTICAST_LOOP (34)
value IP_MULTICAST_TTL (33)
value IP_NODEFRAG (22)
value IP_OPTIONS (4)
value IP_ORIGDSTADDR (20)
value IP_PASSSEC (18)
value IP_PKTINFO (8)
value IP_PKTOPTIONS (9)
value IP_PMTUDISC (10)
value IP_PMTUDISC_DO (2)
value IP_PMTUDISC_DONT (0)
value IP_PMTUDISC_INTERFACE (4)
value IP_PMTUDISC_OMIT (5)
value IP_PMTUDISC_PROBE (3)
value IP_PMTUDISC_WANT (1)
value IP_RECVERR (11)
value IP_RECVFRAGSIZE (25)
value IP_RECVOPTS (6)
value IP_RECVORIGDSTADDR (IP_ORIGDSTADDR)
value IP_RECVRETOPTS (IP_RETOPTS)
value IP_RECVTOS (13)
value IP_RECVTTL (12)
value IP_RETOPTS (7)
value IP_ROUTER_ALERT (5)
value IP_TOS (1)
value IP_TRANSPARENT (19)
value IP_TTL (2)
value IP_UNBLOCK_SOURCE (37)
value IP_UNICAST_IF (50)
value IP_XFRM_POLICY (17)
value ITIMER_PROF (ITIMER_PROF)
value ITIMER_REAL (ITIMER_REAL)
value ITIMER_VIRTUAL (ITIMER_VIRTUAL)
value LITTLE_ENDIAN (__LITTLE_ENDIAN)
value LOCK_EX (2)
value LOCK_NB (4)
value LOCK_SH (1)
value LOCK_UN (8)
value LOGIN_NAME_MAX (256)
value L_INCR (SEEK_CUR)
value L_SET (SEEK_SET)
value L_XTND (SEEK_END)
value MAXNAMLEN (NAME_MAX)
value MAX_CANON (255)
value MAX_INPUT (255)
value MCAST_BLOCK_SOURCE (43)
value MCAST_EXCLUDE (0)
value MCAST_INCLUDE (1)
value MCAST_JOIN_GROUP (42)
value MCAST_JOIN_SOURCE_GROUP (46)
value MCAST_LEAVE_GROUP (45)
value MCAST_LEAVE_SOURCE_GROUP (47)
value MCAST_MSFILTER (48)
value MCAST_UNBLOCK_SOURCE (44)
value MQ_PRIO_MAX (32768)
value MSG_BATCH (MSG_BATCH)
value MSG_CMSG_CLOEXEC (MSG_CMSG_CLOEXEC)
value MSG_CONFIRM (MSG_CONFIRM)
value MSG_CTRUNC (MSG_CTRUNC)
value MSG_DONTROUTE (MSG_DONTROUTE)
value MSG_DONTWAIT (MSG_DONTWAIT)
value MSG_EOR (MSG_EOR)
value MSG_ERRQUEUE (MSG_ERRQUEUE)
value MSG_FASTOPEN (MSG_FASTOPEN)
value MSG_FIN (MSG_FIN)
value MSG_MORE (MSG_MORE)
value MSG_NOSIGNAL (MSG_NOSIGNAL)
value MSG_OOB (MSG_OOB)
value MSG_PEEK (MSG_PEEK)
value MSG_PROXY (MSG_PROXY)
value MSG_RST (MSG_RST)
value MSG_SYN (MSG_SYN)
value MSG_TRUNC (MSG_TRUNC)
value MSG_WAITALL (MSG_WAITALL)
value MSG_WAITFORONE (MSG_WAITFORONE)
value MSG_ZEROCOPY (MSG_ZEROCOPY)
value NAME_MAX (255)
value NETDB_SUCCESS (0)
value NFDBITS (__NFDBITS)
value NGROUPS_MAX (65536)
value NI_DGRAM (16)
value NI_MAXHOST (1025)
value NI_MAXSERV (32)
value NI_NAMEREQD (8)
value NI_NOFQDN (4)
value NI_NUMERICHOST (1)
value NI_NUMERICSERV (2)
value NO_ADDRESS (NO_DATA)
value NO_DATA (4)
value NO_RECOVERY (3)
value O_ACCMODE (0c003)
value O_APPEND (0c2000)
value O_ASYNC (0c20000)
value O_CLOEXEC (__O_CLOEXEC)
value O_CREAT (0c100)
value O_DIRECTORY (__O_DIRECTORY)
value O_DSYNC (__O_DSYNC)
value O_EXCL (0c200)
value O_FSYNC (O_SYNC)
value O_NDELAY (O_NONBLOCK)
value O_NOCTTY (0c400)
value O_NOFOLLOW (__O_NOFOLLOW)
value O_NONBLOCK (0c4000)
value O_RDONLY (00)
value O_RDWR (0c2)
value O_RSYNC (O_SYNC)
value O_SYNC (0c4010000)
value O_TRUNC (0c1000)
value O_WRONLY (0c1)
value PATH_MAX (4096)
value PDP_ENDIAN (__PDP_ENDIAN)
value PF_ALG (38)
value PF_APPLETALK (5)
value PF_ASH (18)
value PF_ATMPVC (8)
value PF_ATMSVC (20)
value PF_BLUETOOTH (31)
value PF_BRIDGE (7)
value PF_CAIF (37)
value PF_CAN (29)
value PF_ECONET (19)
value PF_FILE (PF_LOCAL)
value PF_IB (27)
value PF_INET (2)
value PF_IPX (4)
value PF_IRDA (23)
value PF_ISDN (34)
value PF_IUCV (32)
value PF_KCM (41)
value PF_KEY (15)
value PF_LLC (26)
value PF_LOCAL (1)
value PF_MAX (46)
value PF_MCTP (45)
value PF_MPLS (28)
value PF_NETBEUI (13)
value PF_NETLINK (16)
value PF_NETROM (6)
value PF_NFC (39)
value PF_PACKET (17)
value PF_PHONET (35)
value PF_PPPOX (24)
value PF_QIPCRTR (42)
value PF_RDS (21)
value PF_ROSE (11)
value PF_ROUTE (PF_NETLINK)
value PF_RXRPC (33)
value PF_SECURITY (14)
value PF_SMC (43)
value PF_SNA (22)
value PF_TIPC (30)
value PF_UNIX (PF_LOCAL)
value PF_UNSPEC (0)
value PF_VSOCK (40)
value PF_WANPIPE (25)
value PF_XDP (44)
value PIPE_BUF (4096)
value POSIX_FADV_DONTNEED (__POSIX_FADV_DONTNEED)
value POSIX_FADV_NOREUSE (__POSIX_FADV_NOREUSE)
value POSIX_FADV_NORMAL (0)
value POSIX_FADV_RANDOM (1)
value POSIX_FADV_SEQUENTIAL (2)
value POSIX_FADV_WILLNEED (3)
value PTHREAD_DESTRUCTOR_ITERATIONS (_POSIX_THREAD_DESTRUCTOR_ITERATIONS)
value PTHREAD_KEYS_MAX (1024)
value PTHREAD_STACK_MIN (16384)
value RTSIG_MAX (32)
value R_OK (4)
value SCM_RIGHTS (SCM_RIGHTS)
value SCM_SRCRT (IPV6_RXSRCRT)
value SCM_TIMESTAMP (SO_TIMESTAMP)
value SCM_TIMESTAMPING (SO_TIMESTAMPING)
value SCM_TIMESTAMPING_OPT_STATS (54)
value SCM_TIMESTAMPING_PKTINFO (58)
value SCM_TIMESTAMPNS (SO_TIMESTAMPNS)
value SCM_TXTIME (SO_TXTIME)
value SCM_WIFI_STATUS (SO_WIFI_STATUS)
value SEEK_CUR (1)
value SEEK_END (2)
value SEEK_SET (0)
value SHUT_RD (SHUT_RD)
value SHUT_RDWR (SHUT_RDWR)
value SHUT_WR (SHUT_WR)
value SOCK_CLOEXEC (SOCK_CLOEXEC)
value SOCK_DCCP (SOCK_DCCP)
value SOCK_DGRAM (SOCK_DGRAM)
value SOCK_NONBLOCK (SOCK_NONBLOCK)
value SOCK_PACKET (SOCK_PACKET)
value SOCK_RAW (SOCK_RAW)
value SOCK_RDM (SOCK_RDM)
value SOCK_SEQPACKET (SOCK_SEQPACKET)
value SOCK_STREAM (SOCK_STREAM)
value SOL_AAL (265)
value SOL_ALG (279)
value SOL_ATM (264)
value SOL_BLUETOOTH (274)
value SOL_CAIF (278)
value SOL_DCCP (269)
value SOL_DECNET (261)
value SOL_IP (0)
value SOL_IRDA (266)
value SOL_IUCV (277)
value SOL_KCM (281)
value SOL_LLC (268)
value SOL_NETBEUI (267)
value SOL_NETLINK (270)
value SOL_NFC (280)
value SOL_PACKET (263)
value SOL_PNPIPE (275)
value SOL_RAW (255)
value SOL_RDS (276)
value SOL_RXRPC (272)
value SOL_SOCKET (1)
value SOL_TIPC (271)
value SOL_TLS (282)
value SOL_XDP (283)
value SOMAXCONN (4096)
value SO_ACCEPTCONN (30)
value SO_ATTACH_BPF (50)
value SO_ATTACH_FILTER (26)
value SO_ATTACH_REUSEPORT_CBPF (51)
value SO_ATTACH_REUSEPORT_EBPF (52)
value SO_BINDTODEVICE (25)
value SO_BINDTOIFINDEX (62)
value SO_BPF_EXTENSIONS (48)
value SO_BROADCAST (6)
value SO_BSDCOMPAT (14)
value SO_BUF_LOCK (72)
value SO_BUSY_POLL (46)
value SO_BUSY_POLL_BUDGET (70)
value SO_CNX_ADVICE (53)
value SO_COOKIE (57)
value SO_DEBUG (1)
value SO_DETACH_BPF (SO_DETACH_FILTER)
value SO_DETACH_FILTER (27)
value SO_DETACH_REUSEPORT_BPF (68)
value SO_DOMAIN (39)
value SO_DONTROUTE (5)
value SO_ERROR (4)
value SO_GET_FILTER (SO_ATTACH_FILTER)
value SO_INCOMING_CPU (49)
value SO_INCOMING_NAPI_ID (56)
value SO_KEEPALIVE (9)
value SO_LINGER (13)
value SO_LOCK_FILTER (44)
value SO_MARK (36)
value SO_MAX_PACING_RATE (47)
value SO_MEMINFO (55)
value SO_NETNS_COOKIE (71)
value SO_NOFCS (43)
value SO_NO_CHECK (11)
value SO_OOBINLINE (10)
value SO_PASSCRED (16)
value SO_PASSSEC (34)
value SO_PEEK_OFF (42)
value SO_PEERCRED (17)
value SO_PEERGROUPS (59)
value SO_PEERNAME (28)
value SO_PEERSEC (31)
value SO_PREFER_BUSY_POLL (69)
value SO_PRIORITY (12)
value SO_PROTOCOL (38)
value SO_RCVBUF (8)
value SO_RCVBUFFORCE (33)
value SO_RCVLOWAT (18)
value SO_RCVTIMEO (SO_RCVTIMEO_OLD)
value SO_RCVTIMEO_NEW (66)
value SO_RCVTIMEO_OLD (20)
value SO_REUSEADDR (2)
value SO_REUSEPORT (15)
value SO_RXQ_OVFL (40)
value SO_SECURITY_AUTHENTICATION (22)
value SO_SECURITY_ENCRYPTION_NETWORK (24)
value SO_SECURITY_ENCRYPTION_TRANSPORT (23)
value SO_SELECT_ERR_QUEUE (45)
value SO_SNDBUF (7)
value SO_SNDBUFFORCE (32)
value SO_SNDLOWAT (19)
value SO_SNDTIMEO (SO_SNDTIMEO_OLD)
value SO_SNDTIMEO_NEW (67)
value SO_SNDTIMEO_OLD (21)
value SO_TIMESTAMP (SO_TIMESTAMP_OLD)
value SO_TIMESTAMPING (SO_TIMESTAMPING_OLD)
value SO_TIMESTAMPING_NEW (65)
value SO_TIMESTAMPING_OLD (37)
value SO_TIMESTAMPNS (SO_TIMESTAMPNS_OLD)
value SO_TIMESTAMPNS_NEW (64)
value SO_TIMESTAMPNS_OLD (35)
value SO_TIMESTAMP_NEW (63)
value SO_TIMESTAMP_OLD (29)
value SO_TXTIME (61)
value SO_TYPE (3)
value SO_WIFI_STATUS (41)
value SO_ZEROCOPY (60)
value SSIZE_MAX (LONG_MAX)
value STDERR_FILENO (2)
value STDIN_FILENO (0)
value STDOUT_FILENO (1)
value S_BLKSIZE (512)
value S_IEXEC (S_IXUSR)
value S_IFBLK (__S_IFBLK)
value S_IFCHR (__S_IFCHR)
value S_IFDIR (__S_IFDIR)
value S_IFIFO (__S_IFIFO)
value S_IFLNK (__S_IFLNK)
value S_IFMT (__S_IFMT)
value S_IFREG (__S_IFREG)
value S_IFSOCK (__S_IFSOCK)
value S_IREAD (S_IRUSR)
value S_IRUSR (__S_IREAD)
value S_ISGID (__S_ISGID)
value S_ISUID (__S_ISUID)
value S_ISVTX (__S_ISVTX)
value S_IWRITE (S_IWUSR)
value S_IWUSR (__S_IWRITE)
value S_IXUSR (__S_IEXEC)
value TMP_MAX (238328)
value TRY_AGAIN (2)
value TTY_NAME_MAX (32)
value WCHAR_MAX (__WCHAR_MAX)
value WCHAR_MIN (__WCHAR_MIN)
value W_OK (2)
value XATTR_LIST_MAX (65536)
value XATTR_NAME_MAX (255)
value XATTR_SIZE_MAX (65536)
value X_OK (1)
value _ATFILE_SOURCE (1)
value _BITS_BYTESWAP_H (1)
value _BITS_ENDIANNESS_H (1)
value _BITS_ENDIAN_H (1)
value _BITS_ERRNO_H (1)
value _BITS_POSIX_OPT_H (1)
value _BITS_PTHREADTYPES_ARCH_H (1)
value _BITS_PTHREADTYPES_COMMON_H (1)
value _BITS_SETJMP_H (1)
value _BITS_SOCKADDR_H (1)
value _BITS_STAT_H (1)
value _BITS_STDINT_INTN_H (1)
value _BITS_STDINT_UINTN_H (1)
value _BITS_STDIO_LIM_H (1)
value _BITS_STRUCT_STAT_H (1)
value _BITS_TYPESIZES_H (1)
value _BITS_TYPES_H (1)
value _BITS_UINTN_IDENTITY_H (1)
value _BITS_WCHAR_H (1)
value _CS_GNU_LIBC_VERSION (_CS_GNU_LIBC_VERSION)
value _CS_GNU_LIBPTHREAD_VERSION (_CS_GNU_LIBPTHREAD_VERSION)
value _CS_LFS_CFLAGS (_CS_LFS_CFLAGS)
value _CS_LFS_LDFLAGS (_CS_LFS_LDFLAGS)
value _CS_LFS_LIBS (_CS_LFS_LIBS)
value _CS_LFS_LINTFLAGS (_CS_LFS_LINTFLAGS)
value _CS_PATH (_CS_PATH)
value _DEFAULT_SOURCE (1)
value _DIRENT_H (1)
value _ENDIAN_H (1)
value _ERRNO_H (1)
value _FCNTL_H (1)
value _FEATURES_H (1)
value _GETOPT_CORE_H (1)
value _GETOPT_POSIX_H (1)
value _IOFBF (0)
value _IOLBF (1)
value _IONBF (2)
value _LFS_ASYNCHRONOUS_IO (1)
value _LFS_LARGEFILE (1)
value _NETDB_H (1)
value _NETINET_IN_H (1)
value _PC_ALLOC_SIZE_MIN (_PC_ALLOC_SIZE_MIN)
value _PC_ASYNC_IO (_PC_ASYNC_IO)
value _PC_CHOWN_RESTRICTED (_PC_CHOWN_RESTRICTED)
value _PC_FILESIZEBITS (_PC_FILESIZEBITS)
value _PC_LINK_MAX (_PC_LINK_MAX)
value _PC_MAX_CANON (_PC_MAX_CANON)
value _PC_MAX_INPUT (_PC_MAX_INPUT)
value _PC_NAME_MAX (_PC_NAME_MAX)
value _PC_NO_TRUNC (_PC_NO_TRUNC)
value _PC_PATH_MAX (_PC_PATH_MAX)
value _PC_PIPE_BUF (_PC_PIPE_BUF)
value _PC_PRIO_IO (_PC_PRIO_IO)
value _PC_REC_INCR_XFER_SIZE (_PC_REC_INCR_XFER_SIZE)
value _PC_REC_MAX_XFER_SIZE (_PC_REC_MAX_XFER_SIZE)
value _PC_REC_MIN_XFER_SIZE (_PC_REC_MIN_XFER_SIZE)
value _PC_REC_XFER_ALIGN (_PC_REC_XFER_ALIGN)
value _PC_SOCK_MAXBUF (_PC_SOCK_MAXBUF)
value _PC_SYMLINK_MAX (_PC_SYMLINK_MAX)
value _PC_SYNC_IO (_PC_SYNC_IO)
value _PC_VDISABLE (_PC_VDISABLE)
value _POSIX_ADVISORY_INFO (200809L)
value _POSIX_AIO_LISTIO_MAX (2)
value _POSIX_AIO_MAX (1)
value _POSIX_ARG_MAX (4096)
value _POSIX_ASYNCHRONOUS_IO (200809L)
value _POSIX_ASYNC_IO (1)
value _POSIX_BARRIERS (200809L)
value _POSIX_CHILD_MAX (25)
value _POSIX_CHOWN_RESTRICTED (0)
value _POSIX_CLOCKRES_MIN (20000000)
value _POSIX_CLOCK_SELECTION (200809L)
value _POSIX_CPUTIME (0)
value _POSIX_C_SOURCE (200809L)
value _POSIX_DELAYTIMER_MAX (32)
value _POSIX_FSYNC (200809L)
value _POSIX_HOST_NAME_MAX (255)
value _POSIX_JOB_CONTROL (1)
value _POSIX_LINK_MAX (8)
value _POSIX_LOGIN_NAME_MAX (9)
value _POSIX_MAPPED_FILES (200809L)
value _POSIX_MAX_CANON (255)
value _POSIX_MAX_INPUT (255)
value _POSIX_MEMLOCK (200809L)
value _POSIX_MEMLOCK_RANGE (200809L)
value _POSIX_MEMORY_PROTECTION (200809L)
value _POSIX_MESSAGE_PASSING (200809L)
value _POSIX_MONOTONIC_CLOCK (0)
value _POSIX_MQ_OPEN_MAX (8)
value _POSIX_MQ_PRIO_MAX (32)
value _POSIX_NAME_MAX (14)
value _POSIX_NGROUPS_MAX (8)
value _POSIX_NO_TRUNC (1)
value _POSIX_OPEN_MAX (20)
value _POSIX_PATH_MAX (256)
value _POSIX_PIPE_BUF (512)
value _POSIX_PRIORITIZED_IO (200809L)
value _POSIX_PRIORITY_SCHEDULING (200809L)
value _POSIX_RAW_SOCKETS (200809L)
value _POSIX_READER_WRITER_LOCKS (200809L)
value _POSIX_REALTIME_SIGNALS (200809L)
value _POSIX_REENTRANT_FUNCTIONS (1)
value _POSIX_REGEXP (1)
value _POSIX_RE_DUP_MAX (255)
value _POSIX_RTSIG_MAX (8)
value _POSIX_SAVED_IDS (1)
value _POSIX_SEMAPHORES (200809L)
value _POSIX_SEM_NSEMS_MAX (256)
value _POSIX_SEM_VALUE_MAX (32767)
value _POSIX_SHARED_MEMORY_OBJECTS (200809L)
value _POSIX_SHELL (1)
value _POSIX_SIGQUEUE_MAX (32)
value _POSIX_SOURCE (1)
value _POSIX_SPAWN (200809L)
value _POSIX_SPIN_LOCKS (200809L)
value _POSIX_SSIZE_MAX (32767)
value _POSIX_STREAM_MAX (8)
value _POSIX_SYMLINK_MAX (255)
value _POSIX_SYMLOOP_MAX (8)
value _POSIX_SYNCHRONIZED_IO (200809L)
value _POSIX_THREADS (200809L)
value _POSIX_THREAD_ATTR_STACKADDR (200809L)
value _POSIX_THREAD_ATTR_STACKSIZE (200809L)
value _POSIX_THREAD_CPUTIME (0)
value _POSIX_THREAD_DESTRUCTOR_ITERATIONS (4)
value _POSIX_THREAD_KEYS_MAX (128)
value _POSIX_THREAD_PRIORITY_SCHEDULING (200809L)
value _POSIX_THREAD_PRIO_INHERIT (200809L)
value _POSIX_THREAD_PRIO_PROTECT (200809L)
value _POSIX_THREAD_PROCESS_SHARED (200809L)
value _POSIX_THREAD_ROBUST_PRIO_INHERIT (200809L)
value _POSIX_THREAD_SAFE_FUNCTIONS (200809L)
value _POSIX_THREAD_THREADS_MAX (64)
value _POSIX_TIMEOUTS (200809L)
value _POSIX_TIMERS (200809L)
value _POSIX_TIMER_MAX (32)
value _POSIX_TTY_NAME_MAX (9)
value _POSIX_TZNAME_MAX (6)
value _POSIX_VERSION (200809L)
value _RPC_NETDB_H (1)
value _SC_ADVISORY_INFO (_SC_ADVISORY_INFO)
value _SC_AIO_LISTIO_MAX (_SC_AIO_LISTIO_MAX)
value _SC_AIO_MAX (_SC_AIO_MAX)
value _SC_AIO_PRIO_DELTA_MAX (_SC_AIO_PRIO_DELTA_MAX)
value _SC_ARG_MAX (_SC_ARG_MAX)
value _SC_ASYNCHRONOUS_IO (_SC_ASYNCHRONOUS_IO)
value _SC_ATEXIT_MAX (_SC_ATEXIT_MAX)
value _SC_AVPHYS_PAGES (_SC_AVPHYS_PAGES)
value _SC_BARRIERS (_SC_BARRIERS)
value _SC_BASE (_SC_BASE)
value _SC_BC_BASE_MAX (_SC_BC_BASE_MAX)
value _SC_BC_DIM_MAX (_SC_BC_DIM_MAX)
value _SC_BC_SCALE_MAX (_SC_BC_SCALE_MAX)
value _SC_BC_STRING_MAX (_SC_BC_STRING_MAX)
value _SC_CHARCLASS_NAME_MAX (_SC_CHARCLASS_NAME_MAX)
value _SC_CHAR_BIT (_SC_CHAR_BIT)
value _SC_CHAR_MAX (_SC_CHAR_MAX)
value _SC_CHAR_MIN (_SC_CHAR_MIN)
value _SC_CHILD_MAX (_SC_CHILD_MAX)
value _SC_CLK_TCK (_SC_CLK_TCK)
value _SC_CLOCK_SELECTION (_SC_CLOCK_SELECTION)
value _SC_COLL_WEIGHTS_MAX (_SC_COLL_WEIGHTS_MAX)
value _SC_CPUTIME (_SC_CPUTIME)
value _SC_C_LANG_SUPPORT (_SC_C_LANG_SUPPORT)
value _SC_C_LANG_SUPPORT_R (_SC_C_LANG_SUPPORT_R)
value _SC_DELAYTIMER_MAX (_SC_DELAYTIMER_MAX)
value _SC_DEVICE_IO (_SC_DEVICE_IO)
value _SC_DEVICE_SPECIFIC (_SC_DEVICE_SPECIFIC)
value _SC_DEVICE_SPECIFIC_R (_SC_DEVICE_SPECIFIC_R)
value _SC_EQUIV_CLASS_MAX (_SC_EQUIV_CLASS_MAX)
value _SC_EXPR_NEST_MAX (_SC_EXPR_NEST_MAX)
value _SC_FD_MGMT (_SC_FD_MGMT)
value _SC_FIFO (_SC_FIFO)
value _SC_FILE_ATTRIBUTES (_SC_FILE_ATTRIBUTES)
value _SC_FILE_LOCKING (_SC_FILE_LOCKING)
value _SC_FILE_SYSTEM (_SC_FILE_SYSTEM)
value _SC_FSYNC (_SC_FSYNC)
value _SC_GETGR_R_SIZE_MAX (_SC_GETGR_R_SIZE_MAX)
value _SC_GETPW_R_SIZE_MAX (_SC_GETPW_R_SIZE_MAX)
value _SC_HOST_NAME_MAX (_SC_HOST_NAME_MAX)
value _SC_INT_MAX (_SC_INT_MAX)
value _SC_INT_MIN (_SC_INT_MIN)
value _SC_IOV_MAX (_SC_IOV_MAX)
value _SC_JOB_CONTROL (_SC_JOB_CONTROL)
value _SC_LINE_MAX (_SC_LINE_MAX)
value _SC_LOGIN_NAME_MAX (_SC_LOGIN_NAME_MAX)
value _SC_LONG_BIT (_SC_LONG_BIT)
value _SC_MAPPED_FILES (_SC_MAPPED_FILES)
value _SC_MB_LEN_MAX (_SC_MB_LEN_MAX)
value _SC_MEMLOCK (_SC_MEMLOCK)
value _SC_MEMLOCK_RANGE (_SC_MEMLOCK_RANGE)
value _SC_MEMORY_PROTECTION (_SC_MEMORY_PROTECTION)
value _SC_MESSAGE_PASSING (_SC_MESSAGE_PASSING)
value _SC_MINSIGSTKSZ (_SC_MINSIGSTKSZ)
value _SC_MONOTONIC_CLOCK (_SC_MONOTONIC_CLOCK)
value _SC_MQ_OPEN_MAX (_SC_MQ_OPEN_MAX)
value _SC_MQ_PRIO_MAX (_SC_MQ_PRIO_MAX)
value _SC_MULTI_PROCESS (_SC_MULTI_PROCESS)
value _SC_NETWORKING (_SC_NETWORKING)
value _SC_NGROUPS_MAX (_SC_NGROUPS_MAX)
value _SC_NL_ARGMAX (_SC_NL_ARGMAX)
value _SC_NL_LANGMAX (_SC_NL_LANGMAX)
value _SC_NL_MSGMAX (_SC_NL_MSGMAX)
value _SC_NL_NMAX (_SC_NL_NMAX)
value _SC_NL_SETMAX (_SC_NL_SETMAX)
value _SC_NL_TEXTMAX (_SC_NL_TEXTMAX)
value _SC_NPROCESSORS_CONF (_SC_NPROCESSORS_CONF)
value _SC_NPROCESSORS_ONLN (_SC_NPROCESSORS_ONLN)
value _SC_NZERO (_SC_NZERO)
value _SC_OPEN_MAX (_SC_OPEN_MAX)
value _SC_PAGESIZE (_SC_PAGESIZE)
value _SC_PAGE_SIZE (_SC_PAGESIZE)
value _SC_PASS_MAX (_SC_PASS_MAX)
value _SC_PHYS_PAGES (_SC_PHYS_PAGES)
value _SC_PII (_SC_PII)
value _SC_PII_INTERNET (_SC_PII_INTERNET)
value _SC_PII_INTERNET_DGRAM (_SC_PII_INTERNET_DGRAM)
value _SC_PII_INTERNET_STREAM (_SC_PII_INTERNET_STREAM)
value _SC_PII_OSI (_SC_PII_OSI)
value _SC_PII_OSI_CLTS (_SC_PII_OSI_CLTS)
value _SC_PII_OSI_COTS (_SC_PII_OSI_COTS)
value _SC_PII_OSI_M (_SC_PII_OSI_M)
value _SC_PII_SOCKET (_SC_PII_SOCKET)
value _SC_PII_XTI (_SC_PII_XTI)
value _SC_PIPE (_SC_PIPE)
value _SC_POLL (_SC_POLL)
value _SC_PRIORITIZED_IO (_SC_PRIORITIZED_IO)
value _SC_PRIORITY_SCHEDULING (_SC_PRIORITY_SCHEDULING)
value _SC_RAW_SOCKETS (_SC_RAW_SOCKETS)
value _SC_READER_WRITER_LOCKS (_SC_READER_WRITER_LOCKS)
value _SC_REALTIME_SIGNALS (_SC_REALTIME_SIGNALS)
value _SC_REGEXP (_SC_REGEXP)
value _SC_REGEX_VERSION (_SC_REGEX_VERSION)
value _SC_RE_DUP_MAX (_SC_RE_DUP_MAX)
value _SC_RTSIG_MAX (_SC_RTSIG_MAX)
value _SC_SAVED_IDS (_SC_SAVED_IDS)
value _SC_SCHAR_MAX (_SC_SCHAR_MAX)
value _SC_SCHAR_MIN (_SC_SCHAR_MIN)
value _SC_SELECT (_SC_SELECT)
value _SC_SEMAPHORES (_SC_SEMAPHORES)
value _SC_SEM_NSEMS_MAX (_SC_SEM_NSEMS_MAX)
value _SC_SEM_VALUE_MAX (_SC_SEM_VALUE_MAX)
value _SC_SHARED_MEMORY_OBJECTS (_SC_SHARED_MEMORY_OBJECTS)
value _SC_SHELL (_SC_SHELL)
value _SC_SHRT_MAX (_SC_SHRT_MAX)
value _SC_SHRT_MIN (_SC_SHRT_MIN)
value _SC_SIGNALS (_SC_SIGNALS)
value _SC_SIGQUEUE_MAX (_SC_SIGQUEUE_MAX)
value _SC_SIGSTKSZ (_SC_SIGSTKSZ)
value _SC_SINGLE_PROCESS (_SC_SINGLE_PROCESS)
value _SC_SPAWN (_SC_SPAWN)
value _SC_SPIN_LOCKS (_SC_SPIN_LOCKS)
value _SC_SPORADIC_SERVER (_SC_SPORADIC_SERVER)
value _SC_SSIZE_MAX (_SC_SSIZE_MAX)
value _SC_SS_REPL_MAX (_SC_SS_REPL_MAX)
value _SC_STREAMS (_SC_STREAMS)
value _SC_STREAM_MAX (_SC_STREAM_MAX)
value _SC_SYMLOOP_MAX (_SC_SYMLOOP_MAX)
value _SC_SYNCHRONIZED_IO (_SC_SYNCHRONIZED_IO)
value _SC_SYSTEM_DATABASE (_SC_SYSTEM_DATABASE)
value _SC_SYSTEM_DATABASE_R (_SC_SYSTEM_DATABASE_R)
value _SC_THREADS (_SC_THREADS)
value _SC_THREAD_ATTR_STACKADDR (_SC_THREAD_ATTR_STACKADDR)
value _SC_THREAD_ATTR_STACKSIZE (_SC_THREAD_ATTR_STACKSIZE)
value _SC_THREAD_CPUTIME (_SC_THREAD_CPUTIME)
value _SC_THREAD_DESTRUCTOR_ITERATIONS (_SC_THREAD_DESTRUCTOR_ITERATIONS)
value _SC_THREAD_KEYS_MAX (_SC_THREAD_KEYS_MAX)
value _SC_THREAD_PRIORITY_SCHEDULING (_SC_THREAD_PRIORITY_SCHEDULING)
value _SC_THREAD_PRIO_INHERIT (_SC_THREAD_PRIO_INHERIT)
value _SC_THREAD_PRIO_PROTECT (_SC_THREAD_PRIO_PROTECT)
value _SC_THREAD_PROCESS_SHARED (_SC_THREAD_PROCESS_SHARED)
value _SC_THREAD_ROBUST_PRIO_INHERIT (_SC_THREAD_ROBUST_PRIO_INHERIT)
value _SC_THREAD_ROBUST_PRIO_PROTECT (_SC_THREAD_ROBUST_PRIO_PROTECT)
value _SC_THREAD_SAFE_FUNCTIONS (_SC_THREAD_SAFE_FUNCTIONS)
value _SC_THREAD_SPORADIC_SERVER (_SC_THREAD_SPORADIC_SERVER)
value _SC_THREAD_STACK_MIN (_SC_THREAD_STACK_MIN)
value _SC_THREAD_THREADS_MAX (_SC_THREAD_THREADS_MAX)
value _SC_TIMEOUTS (_SC_TIMEOUTS)
value _SC_TIMERS (_SC_TIMERS)
value _SC_TIMER_MAX (_SC_TIMER_MAX)
value _SC_TRACE (_SC_TRACE)
value _SC_TRACE_EVENT_FILTER (_SC_TRACE_EVENT_FILTER)
value _SC_TRACE_EVENT_NAME_MAX (_SC_TRACE_EVENT_NAME_MAX)
value _SC_TRACE_INHERIT (_SC_TRACE_INHERIT)
value _SC_TRACE_LOG (_SC_TRACE_LOG)
value _SC_TRACE_NAME_MAX (_SC_TRACE_NAME_MAX)
value _SC_TRACE_SYS_MAX (_SC_TRACE_SYS_MAX)
value _SC_TRACE_USER_EVENT_MAX (_SC_TRACE_USER_EVENT_MAX)
value _SC_TTY_NAME_MAX (_SC_TTY_NAME_MAX)
value _SC_TYPED_MEMORY_OBJECTS (_SC_TYPED_MEMORY_OBJECTS)
value _SC_TZNAME_MAX (_SC_TZNAME_MAX)
value _SC_T_IOV_MAX (_SC_T_IOV_MAX)
value _SC_UCHAR_MAX (_SC_UCHAR_MAX)
value _SC_UINT_MAX (_SC_UINT_MAX)
value _SC_UIO_MAXIOV (_SC_UIO_MAXIOV)
value _SC_ULONG_MAX (_SC_ULONG_MAX)
value _SC_USER_GROUPS (_SC_USER_GROUPS)
value _SC_USER_GROUPS_R (_SC_USER_GROUPS_R)
value _SC_USHRT_MAX (_SC_USHRT_MAX)
value _SC_VERSION (_SC_VERSION)
value _SC_WORD_BIT (_SC_WORD_BIT)
value _SC_XOPEN_CRYPT (_SC_XOPEN_CRYPT)
value _SC_XOPEN_LEGACY (_SC_XOPEN_LEGACY)
value _SC_XOPEN_REALTIME (_SC_XOPEN_REALTIME)
value _SC_XOPEN_REALTIME_THREADS (_SC_XOPEN_REALTIME_THREADS)
value _SC_XOPEN_SHM (_SC_XOPEN_SHM)
value _SC_XOPEN_STREAMS (_SC_XOPEN_STREAMS)
value _SC_XOPEN_UNIX (_SC_XOPEN_UNIX)
value _SC_XOPEN_VERSION (_SC_XOPEN_VERSION)
value _SC_XOPEN_XCU_VERSION (_SC_XOPEN_XCU_VERSION)
value _SETJMP_H (1)
value _SS_SIZE (128)
value _STDC_PREDEF_H (1)
value _STDINT_H (1)
value _STDIO_H (1)
value _STRUCT_TIMESPEC (1)
value _SYS_CDEFS_H (1)
value _SYS_EPOLL_H (1)
value _SYS_POLL_H (1)
value _SYS_SELECT_H (1)
value _SYS_SOCKET_H (1)
value _SYS_STAT_H (1)
value _SYS_TIME_H (1)
value _SYS_TYPES_H (1)
value _THREAD_MUTEX_INTERNAL_H (1)
value _THREAD_SHARED_TYPES_H (1)
value _UNISTD_H (1)
value _XOPEN_LEGACY (1)
value _XOPEN_REALTIME (1)
value _XOPEN_REALTIME_THREADS (1)
value _XOPEN_SHM (1)
value _XOPEN_UNIX (1)
value _XOPEN_VERSION (700)
value _XOPEN_XCU_VERSION (4)
value __ATOMIC_ACQUIRE (2)
value __ATOMIC_ACQ_REL (4)
value __ATOMIC_CONSUME (1)
value __ATOMIC_RELAXED (0)
value __ATOMIC_RELEASE (3)
value __ATOMIC_SEQ_CST (5)
value __BIGGEST_ALIGNMENT__ (16)
value __BIG_ENDIAN (4321)
value __BITINT_MAXWIDTH__ (128)
value __BITS_PER_LONG (64)
value __BIT_TYPES_DEFINED__ (1)
value __BLKCNT_T_TYPE (__SYSCALL_SLONG_TYPE)
value __BLKSIZE_T_TYPE (__SYSCALL_SLONG_TYPE)
value __BOOL_WIDTH__ (8)
value __BYTE_ORDER (__LITTLE_ENDIAN)
value __BYTE_ORDER__ (__ORDER_LITTLE_ENDIAN__)
value __CHAR_BIT__ (8)
value __CLANG_ATOMIC_BOOL_LOCK_FREE (2)
value __CLANG_ATOMIC_CHAR_LOCK_FREE (2)
value __CLANG_ATOMIC_INT_LOCK_FREE (2)
value __CLANG_ATOMIC_LLONG_LOCK_FREE (2)
value __CLANG_ATOMIC_LONG_LOCK_FREE (2)
value __CLANG_ATOMIC_POINTER_LOCK_FREE (2)
value __CLANG_ATOMIC_SHORT_LOCK_FREE (2)
value __CLANG_ATOMIC_WCHAR_T_LOCK_FREE (2)
value __CLOCKID_T_TYPE (__S32_TYPE)
value __CLOCK_T_TYPE (__SYSCALL_SLONG_TYPE)
value __CONSTANT_CFSTRINGS__ (1)
value __CPU_MASK_TYPE (__SYSCALL_ULONG_TYPE)
value __DADDR_T_TYPE (__S32_TYPE)
value __DBL_DECIMAL_DIG__ (17)
value __DBL_DIG__ (15)
value __DBL_HAS_DENORM__ (1)
value __DBL_HAS_INFINITY__ (1)
value __DBL_HAS_QUIET_NAN__ (1)
value __DBL_MANT_DIG__ (53)
value __DBL_MAX_EXP__ (1024)
value __DECIMAL_DIG__ (__LDBL_DECIMAL_DIG__)
value __DEV_T_TYPE (__UQUAD_TYPE)
value __ELF__ (1)
value __FD_SETSIZE (1024)
value __FINITE_MATH_ONLY__ (0)
value __FLOAT_WORD_ORDER (__BYTE_ORDER)
value __FLT_DECIMAL_DIG__ (9)
value __FLT_DIG__ (6)
value __FLT_HAS_DENORM__ (1)
value __FLT_HAS_INFINITY__ (1)
value __FLT_HAS_QUIET_NAN__ (1)
value __FLT_MANT_DIG__ (24)
value __FLT_MAX_EXP__ (128)
value __FLT_RADIX__ (2)
value __FSBLKCNT_T_TYPE (__SYSCALL_ULONG_TYPE)
value __FSFILCNT_T_TYPE (__SYSCALL_ULONG_TYPE)
value __FSWORD_T_TYPE (__SYSCALL_SLONG_TYPE)
value __FXSR__ (1)
value __F_GETOWN (9)
value __F_GETOWN_EX (16)
value __F_GETSIG (11)
value __F_SETOWN (8)
value __F_SETOWN_EX (15)
value __F_SETSIG (10)
value __GCC_ASM_FLAG_OUTPUTS__ (1)
value __GCC_ATOMIC_BOOL_LOCK_FREE (2)
value __GCC_ATOMIC_CHAR_LOCK_FREE (2)
value __GCC_ATOMIC_INT_LOCK_FREE (2)
value __GCC_ATOMIC_LLONG_LOCK_FREE (2)
value __GCC_ATOMIC_LONG_LOCK_FREE (2)
value __GCC_ATOMIC_POINTER_LOCK_FREE (2)
value __GCC_ATOMIC_SHORT_LOCK_FREE (2)
value __GCC_ATOMIC_TEST_AND_SET_TRUEVAL (1)
value __GCC_ATOMIC_WCHAR_T_LOCK_FREE (2)
value __GID_T_TYPE (__U32_TYPE)
value __GLIBC_MINOR__ (35)
value __GLIBC_USE_DEPRECATED_GETS (0)
value __GLIBC_USE_DEPRECATED_SCANF (0)
value __GLIBC__ (2)
value __GNUC_MINOR__ (2)
value __GNUC_PATCHLEVEL__ (1)
value __GNUC_STDC_INLINE__ (1)
value __GNUC_VA_LIST (1)
value __GNUC__ (4)
value __GNU_LIBRARY__ (6)
value __GXX_ABI_VERSION (1002)
value __HAVE_FLOATN_NOT_TYPEDEF (0)
value __HAVE_GENERIC_SELECTION (1)
value __ID_T_TYPE (__U32_TYPE)
value __INO_T_TYPE (__SYSCALL_ULONG_TYPE)
value __INTMAX_C_SUFFIX__ (L)
value __INTMAX_MAX__ (9223372036854775807L)
value __INTMAX_WIDTH__ (64)
value __INTPTR_MAX__ (9223372036854775807L)
value __INTPTR_WIDTH__ (64)
value __INT_MAX__ (2147483647)
value __INT_WIDTH__ (32)
value __KEY_T_TYPE (__S32_TYPE)
value __LDBL_DECIMAL_DIG__ (21)
value __LDBL_DIG__ (18)
value __LDBL_HAS_DENORM__ (1)
value __LDBL_HAS_INFINITY__ (1)
value __LDBL_HAS_QUIET_NAN__ (1)
value __LDBL_MANT_DIG__ (64)
value __LDBL_MAX_EXP__ (16384)
value __LITTLE_ENDIAN (1234)
value __LITTLE_ENDIAN__ (1)
value __LLONG_WIDTH__ (64)
value __LONG_LONG_MAX__ (9223372036854775807LL)
value __LONG_MAX__ (9223372036854775807L)
value __LONG_WIDTH__ (64)
value __MMX__ (1)
value __MODE_T_TYPE (__U32_TYPE)
value __NLINK_T_TYPE (__SYSCALL_ULONG_TYPE)
value __NO_INLINE__ (1)
value __NO_MATH_INLINES (1)
value __OBJC_BOOL_IS_BOOL (0)
value __OFF_T_TYPE (__SYSCALL_SLONG_TYPE)
value __OPENCL_MEMORY_SCOPE_ALL_SVM_DEVICES (3)
value __OPENCL_MEMORY_SCOPE_DEVICE (2)
value __OPENCL_MEMORY_SCOPE_SUB_GROUP (4)
value __OPENCL_MEMORY_SCOPE_WORK_GROUP (1)
value __OPENCL_MEMORY_SCOPE_WORK_ITEM (0)
value __ORDER_BIG_ENDIAN__ (4321)
value __ORDER_LITTLE_ENDIAN__ (1234)
value __ORDER_PDP_ENDIAN__ (3412)
value __O_CLOEXEC (0c2000000)
value __O_DIRECT (0c40000)
value __O_DIRECTORY (0c200000)
value __O_DSYNC (0c10000)
value __O_LARGEFILE (0)
value __O_NOATIME (0c1000000)
value __O_NOFOLLOW (0c400000)
value __O_PATH (0c10000000)
value __PDP_ENDIAN (3412)
value __PIC__ (2)
value __PID_T_TYPE (__S32_TYPE)
value __PIE__ (2)
value __POINTER_WIDTH__ (64)
value __POSIX_FADV_DONTNEED (4)
value __POSIX_FADV_NOREUSE (5)
value __PRAGMA_REDEFINE_EXTNAME (1)
value __PTHREAD_MUTEX_HAVE_PREV (1)
value __PTRDIFF_MAX__ (9223372036854775807L)
value __PTRDIFF_WIDTH__ (64)
value __RLIM_T_TYPE (__SYSCALL_ULONG_TYPE)
value __SCHAR_MAX__ (127)
value __SEG_FS (1)
value __SEG_GS (1)
value __SHRT_MAX__ (32767)
value __SHRT_WIDTH__ (16)
value __SIG_ATOMIC_MAX__ (2147483647)
value __SIG_ATOMIC_WIDTH__ (32)
value __SIZEOF_DOUBLE__ (8)
value __SIZEOF_FLOAT__ (4)
value __SIZEOF_INT__ (4)
value __SIZEOF_LONG_DOUBLE__ (16)
value __SIZEOF_LONG_LONG__ (8)
value __SIZEOF_LONG__ (8)
value __SIZEOF_POINTER__ (8)
value __SIZEOF_PTHREAD_ATTR_T (56)
value __SIZEOF_PTHREAD_BARRIERATTR_T (4)
value __SIZEOF_PTHREAD_BARRIER_T (32)
value __SIZEOF_PTHREAD_CONDATTR_T (4)
value __SIZEOF_PTHREAD_COND_T (48)
value __SIZEOF_PTHREAD_MUTEXATTR_T (4)
value __SIZEOF_PTHREAD_MUTEX_T (40)
value __SIZEOF_PTHREAD_RWLOCKATTR_T (8)
value __SIZEOF_PTHREAD_RWLOCK_T (56)
value __SIZEOF_PTRDIFF_T__ (8)
value __SIZEOF_SHORT__ (2)
value __SIZEOF_SIZE_T__ (8)
value __SIZEOF_WCHAR_T__ (4)
value __SIZEOF_WINT_T__ (4)
value __SIZE_MAX__ (18446744073709551615UL)
value __SIZE_WIDTH__ (64)
value __SSE_MATH__ (1)
value __SSE__ (1)
value __SSIZE_T_TYPE (__SWORD_TYPE)
value __STDC_HOSTED__ (1)
value __STDC_VERSION__ (201710L)
value __STDC__ (1)
value __SUSECONDS_T_TYPE (__SYSCALL_SLONG_TYPE)
value __SYSCALL_SLONG_TYPE (__SLONGWORD_TYPE)
value __SYSCALL_ULONG_TYPE (__ULONGWORD_TYPE)
value __SYSCALL_WORDSIZE (64)
value __S_IEXEC (0c100)
value __S_IFBLK (0c060000)
value __S_IFCHR (0c020000)
value __S_IFDIR (0c040000)
value __S_IFIFO (0c010000)
value __S_IFLNK (0c120000)
value __S_IFMT (0c170000)
value __S_IFREG (0c100000)
value __S_IFSOCK (0c140000)
value __S_IREAD (0c400)
value __S_ISGID (0c2000)
value __S_ISUID (0c4000)
value __S_ISVTX (0c1000)
value __S_IWRITE (0c200)
value __TIMESIZE (__WORDSIZE)
value __TIME_T_TYPE (__SYSCALL_SLONG_TYPE)
value __UID_T_TYPE (__U32_TYPE)
value __UINTMAX_C_SUFFIX__ (UL)
value __UINTMAX_MAX__ (18446744073709551615UL)
value __UINTMAX_WIDTH__ (64)
value __UINTPTR_MAX__ (18446744073709551615UL)
value __UINTPTR_WIDTH__ (64)
value __USECONDS_T_TYPE (__U32_TYPE)
value __USE_ATFILE (1)
value __USE_FORTIFY_LEVEL (0)
value __USE_MISC (1)
value __USE_POSIX (1)
value __USE_POSIX_IMPLICITLY (1)
value __WCHAR_MAX (__WCHAR_MAX__)
value __WCHAR_MAX__ (2147483647)
value __WCHAR_WIDTH__ (32)
value __WINT_MAX__ (4294967295U)
value __WINT_UNSIGNED__ (1)
value __WINT_WIDTH__ (32)
value __WORDSIZE (64)

