
value EAGAIN (35)
value SOCK_STREAM (1)
value F_GETFL (3)
value F_SETFL (4)
value O_NONBLOCK (4)

value SOL_SOCKET (65535)
value SO_REUSEADDR (4)
value SO_RCVTIMEO (4102)

value AF_INET (2)
value AF_UNIX (1)

value AI_PASSIVE (1)
value AI_CANONNAME (2)
value AI_NUMERICHOST (4)

value POLLIN (1)
value POLLOUT (4)
value POLLERR (8)
value POLLHUP (16)
value POLLRDHUP (8192)
