
value ACCESSX_MAX_DESCRIPTORS (100)
value AF_APPLETALK (16)
value AF_CCITT (10)
value AF_CHAOS (5)
value AF_CNT (21)
value AF_COIP (20)
value AF_DATAKIT (9)
value AF_DLI (13)
value AF_ECMA (8)
value AF_HYLINK (15)
value AF_IMPLINK (3)
value AF_INET (2)
value AF_IPX (23)
value AF_ISDN (28)
value AF_ISO (7)
value AF_LAT (14)
value AF_LINK (18)
value AF_LOCAL (AF_UNIX)
value AF_MAX (41)
value AF_NATM (31)
value AF_NDRV (27)
value AF_NETBIOS (33)
value AF_NS (6)
value AF_OSI (AF_ISO)
value AF_PPP (34)
value AF_PUP (4)
value AF_ROUTE (17)
value AF_SIP (24)
value AF_SNA (11)
value AF_SYSTEM (32)
value AF_UNIX (1)
value AF_UNSPEC (0)
value AF_UTUN (38)
value AF_VSOCK (40)
value BADSIG (SIG_ERR)
value BIG_ENDIAN (__DARWIN_BIG_ENDIAN)
value BUFSIZ (1024)
value BUS_ADRALN (1)
value BUS_ADRERR (2)
value BUS_NOOP (0)
value BUS_OBJERR (3)
value BYTE_ORDER (__DARWIN_BYTE_ORDER)
value CLD_CONTINUED (6)
value CLD_DUMPED (3)
value CLD_EXITED (1)
value CLD_KILLED (2)
value CLD_NOOP (0)
value CLD_STOPPED (5)
value CLD_TRAPPED (4)
value CLOCKS_PER_SEC (1000000)
value CLOCK_MONOTONIC (_CLOCK_MONOTONIC)
value CLOCK_MONOTONIC_RAW (_CLOCK_MONOTONIC_RAW)
value CLOCK_MONOTONIC_RAW_APPROX (_CLOCK_MONOTONIC_RAW_APPROX)
value CLOCK_PROCESS_CPUTIME_ID (_CLOCK_PROCESS_CPUTIME_ID)
value CLOCK_REALTIME (_CLOCK_REALTIME)
value CLOCK_THREAD_CPUTIME_ID (_CLOCK_THREAD_CPUTIME_ID)
value CLOCK_UPTIME_RAW (_CLOCK_UPTIME_RAW)
value CLOCK_UPTIME_RAW_APPROX (_CLOCK_UPTIME_RAW_APPROX)
value DIRBLKSIZ (1024)
value DST_AUST (2)
value DST_CAN (6)
value DST_EET (5)
value DST_MET (4)
value DST_NONE (0)
value DST_USA (1)
value DST_WET (3)
value DT_BLK (6)
value DT_CHR (2)
value DT_DIR (4)
value DT_FIFO (1)
value DT_LNK (10)
value DT_REG (8)
value DT_SOCK (12)
value DT_UNKNOWN (0)
value DT_WHT (14)
value EACCES (13)
value EADDRINUSE (48)
value EADDRNOTAVAIL (49)
value EAFNOSUPPORT (47)
value EAGAIN (35)
value EAI_ADDRFAMILY (1)
value EAI_AGAIN (2)
value EAI_BADFLAGS (3)
value EAI_BADHINTS (12)
value EAI_FAIL (4)
value EAI_FAMILY (5)
value EAI_MAX (15)
value EAI_MEMORY (6)
value EAI_NODATA (7)
value EAI_NONAME (8)
value EAI_OVERFLOW (14)
value EAI_PROTOCOL (13)
value EAI_SERVICE (9)
value EAI_SOCKTYPE (10)
value EAI_SYSTEM (11)
value EALREADY (37)
value EAUTH (80)
value EBADARCH (86)
value EBADEXEC (85)
value EBADF (9)
value EBADMACHO (88)
value EBADMSG (94)
value EBADRPC (72)
value EBUSY (16)
value ECANCELED (89)
value ECHILD (10)
value ECONNABORTED (53)
value ECONNREFUSED (61)
value ECONNRESET (54)
value EDEADLK (11)
value EDESTADDRREQ (39)
value EDEVERR (83)
value EDOM (33)
value EDQUOT (69)
value EEXIST (17)
value EFAULT (14)
value EFBIG (27)
value EFTYPE (79)
value EHOSTDOWN (64)
value EHOSTUNREACH (65)
value EIDRM (90)
value EILSEQ (92)
value EINPROGRESS (36)
value EINTR (4)
value EINVAL (22)
value EIO (5)
value EISCONN (56)
value EISDIR (21)
value ELAST (106)
value ELOOP (62)
value EMFILE (24)
value EMLINK (31)
value EMSGSIZE (40)
value EMULTIHOP (95)
value ENAMETOOLONG (63)
value ENEEDAUTH (81)
value ENETDOWN (50)
value ENETRESET (52)
value ENETUNREACH (51)
value ENFILE (23)
value ENOATTR (93)
value ENOBUFS (55)
value ENODATA (96)
value ENODEV (19)
value ENOENT (2)
value ENOEXEC (8)
value ENOLCK (77)
value ENOLINK (97)
value ENOMEM (12)
value ENOMSG (91)
value ENOPOLICY (103)
value ENOPROTOOPT (42)
value ENOSPC (28)
value ENOSR (98)
value ENOSTR (99)
value ENOSYS (78)
value ENOTBLK (15)
value ENOTCONN (57)
value ENOTDIR (20)
value ENOTEMPTY (66)
value ENOTRECOVERABLE (104)
value ENOTSOCK (38)
value ENOTSUP (45)
value ENOTTY (25)
value ENXIO (6)
value EOPNOTSUPP (102)
value EOVERFLOW (84)
value EOWNERDEAD (105)
value EPERM (1)
value EPFNOSUPPORT (46)
value EPIPE (32)
value EPROCLIM (67)
value EPROCUNAVAIL (76)
value EPROGMISMATCH (75)
value EPROGUNAVAIL (74)
value EPROTO (100)
value EPROTONOSUPPORT (43)
value EPROTOTYPE (41)
value EPWROFF (82)
value EQFULL (106)
value ERANGE (34)
value EREMOTE (71)
value EROFS (30)
value ERPCMISMATCH (73)
value ESHLIBVERS (87)
value ESHUTDOWN (58)
value ESOCKTNOSUPPORT (44)
value ESPIPE (29)
value ESRCH (3)
value ESTALE (70)
value ETIME (101)
value ETIMEDOUT (60)
value ETOOMANYREFS (59)
value ETXTBSY (26)
value EUSERS (68)
value EWOULDBLOCK (EAGAIN)
value EXDEV (18)
value EXIT_FAILURE (1)
value EXIT_SUCCESS (0)
value FAPPEND (O_APPEND)
value FASYNC (O_ASYNC)
value FD_CLOEXEC (1)
value FD_SETSIZE (__DARWIN_FD_SETSIZE)
value FFDSYNC (O_DSYNC)
value FFSYNC (O_FSYNC)
value FILENAME_MAX (1024)
value FILESEC_GUID (FILESEC_UUID)
value FNDELAY (O_NONBLOCK)
value FNONBLOCK (O_NONBLOCK)
value FOPEN_MAX (20)
value FPE_FLTDIV (1)
value FPE_FLTINV (5)
value FPE_FLTOVF (2)
value FPE_FLTRES (4)
value FPE_FLTSUB (6)
value FPE_FLTUND (3)
value FPE_INTDIV (7)
value FPE_INTOVF (8)
value FPE_NOOP (0)
value F_ADDFILESIGS (61)
value F_ADDFILESIGS_FOR_DYLD_SIM (83)
value F_ADDFILESIGS_INFO (103)
value F_ADDFILESIGS_RETURN (97)
value F_ADDFILESUPPL (104)
value F_ADDSIGS (59)
value F_BARRIERFSYNC (85)
value F_CHECK_LV (98)
value F_CHKCLEAN (41)
value F_DUPFD (0)
value F_DUPFD_CLOEXEC (67)
value F_FINDSIGS (78)
value F_FLUSH_DATA (40)
value F_FREEZE_FS (53)
value F_FULLFSYNC (51)
value F_GETCODEDIR (72)
value F_GETFD (1)
value F_GETFL (3)
value F_GETLK (7)
value F_GETLKPID (66)
value F_GETNOSIGPIPE (74)
value F_GETOWN (5)
value F_GETPATH (50)
value F_GETPATH_MTMINFO (71)
value F_GETPATH_NOFIRMLINK (102)
value F_GETPROTECTIONCLASS (63)
value F_GETPROTECTIONLEVEL (77)
value F_GETSIGSINFO (105)
value F_GLOBAL_NOCACHE (55)
value F_LOCK (1)
value F_NOCACHE (48)
value F_NODIRECT (62)
value F_OK (0)
value F_PATHPKG_CHECK (52)
value F_PEOFPOSMODE (3)
value F_PREALLOCATE (42)
value F_PUNCHHOLE (99)
value F_RDADVISE (44)
value F_RDAHEAD (45)
value F_RDLCK (1)
value F_SETBACKINGSTORE (70)
value F_SETFD (2)
value F_SETFL (4)
value F_SETLK (8)
value F_SETLKW (9)
value F_SETLKWTIMEOUT (10)
value F_SETNOSIGPIPE (73)
value F_SETOWN (6)
value F_SETPROTECTIONCLASS (64)
value F_SETSIZE (43)
value F_SINGLE_WRITER (76)
value F_SPECULATIVE_READ (101)
value F_TEST (3)
value F_THAW_FS (54)
value F_TLOCK (2)
value F_TRANSCODEKEY (75)
value F_TRIM_ACTIVE_FILE (100)
value F_ULOCK (0)
value F_UNLCK (2)
value F_VOLPOSMODE (4)
value F_WRLCK (3)
value GETSIGSINFO_PLATFORM_BINARY (1)
value HOST_NOT_FOUND (1)
value ILL_BADSTK (8)
value ILL_COPROC (7)
value ILL_ILLADR (5)
value ILL_ILLOPC (1)
value ILL_ILLOPN (4)
value ILL_ILLTRP (2)
value ILL_NOOP (0)
value ILL_PRVOPC (3)
value ILL_PRVREG (6)
value INET_ADDRSTRLEN (16)
value INTPTR_MAX (9223372036854775807L)
value IN_CLASSA_MAX (128)
value IN_CLASSA_NSHIFT (24)
value IN_CLASSB_MAX (65536)
value IN_CLASSB_NSHIFT (16)
value IN_CLASSC_NSHIFT (8)
value IN_CLASSD_NSHIFT (28)
value IN_LOOPBACKNET (127)
value IOPOL_APPLICATION (IOPOL_STANDARD)
value IOPOL_ATIME_UPDATES_DEFAULT (0)
value IOPOL_ATIME_UPDATES_OFF (1)
value IOPOL_DEFAULT (0)
value IOPOL_IMPORTANT (1)
value IOPOL_MATERIALIZE_DATALESS_FILES_DEFAULT (0)
value IOPOL_MATERIALIZE_DATALESS_FILES_OFF (1)
value IOPOL_MATERIALIZE_DATALESS_FILES_ON (2)
value IOPOL_NORMAL (IOPOL_IMPORTANT)
value IOPOL_PASSIVE (2)
value IOPOL_SCOPE_DARWIN_BG (2)
value IOPOL_SCOPE_PROCESS (0)
value IOPOL_SCOPE_THREAD (1)
value IOPOL_STANDARD (5)
value IOPOL_THROTTLE (3)
value IOPOL_TYPE_DISK (0)
value IOPOL_TYPE_VFS_ATIME_UPDATES (2)
value IOPOL_TYPE_VFS_IGNORE_CONTENT_PROTECTION (6)
value IOPOL_TYPE_VFS_IGNORE_PERMISSIONS (7)
value IOPOL_TYPE_VFS_MATERIALIZE_DATALESS_FILES (3)
value IOPOL_TYPE_VFS_SKIP_MTIME_UPDATE (8)
value IOPOL_TYPE_VFS_STATFS_NO_DATA_VOLUME (4)
value IOPOL_TYPE_VFS_TRIGGER_RESOLVE (5)
value IOPOL_UTILITY (4)
value IOPOL_VFS_CONTENT_PROTECTION_DEFAULT (0)
value IOPOL_VFS_CONTENT_PROTECTION_IGNORE (1)
value IOPOL_VFS_IGNORE_PERMISSIONS_OFF (0)
value IOPOL_VFS_IGNORE_PERMISSIONS_ON (1)
value IOPOL_VFS_SKIP_MTIME_UPDATE_OFF (0)
value IOPOL_VFS_SKIP_MTIME_UPDATE_ON (1)
value IOPOL_VFS_STATFS_FORCE_NO_DATA_VOLUME (1)
value IOPOL_VFS_STATFS_NO_DATA_VOLUME_DEFAULT (0)
value IOPOL_VFS_TRIGGER_RESOLVE_DEFAULT (0)
value IOPOL_VFS_TRIGGER_RESOLVE_OFF (1)
value IPCTL_ACCEPTSOURCEROUTE (13)
value IPCTL_DEFTTL (3)
value IPCTL_DIRECTEDBROADCAST (9)
value IPCTL_FASTFORWARDING (14)
value IPCTL_FORWARDING (1)
value IPCTL_GIF_TTL (16)
value IPCTL_INTRQDROPS (11)
value IPCTL_INTRQMAXLEN (10)
value IPCTL_KEEPFAITH (15)
value IPCTL_MAXID (17)
value IPCTL_RTEXPIRE (5)
value IPCTL_RTMAXCACHE (7)
value IPCTL_RTMINEXPIRE (6)
value IPCTL_SENDREDIRECTS (2)
value IPCTL_SOURCEROUTE (8)
value IPCTL_STATS (12)
value IPPORT_HIFIRSTAUTO (49152)
value IPPORT_HILASTAUTO (65535)
value IPPORT_RESERVED (__DARWIN_IPPORT_RESERVED)
value IPPORT_RESERVEDSTART (600)
value IPPORT_USERRESERVED (5000)
value IPPROTO_ADFS (68)
value IPPROTO_AH (51)
value IPPROTO_AHIP (61)
value IPPROTO_APES (99)
value IPPROTO_ARGUS (13)
value IPPROTO_BHA (49)
value IPPROTO_BLT (30)
value IPPROTO_BRSATMON (76)
value IPPROTO_CFTP (62)
value IPPROTO_CHAOS (16)
value IPPROTO_CMTP (38)
value IPPROTO_CPHB (73)
value IPPROTO_CPNX (72)
value IPPROTO_DDP (37)
value IPPROTO_DGP (86)
value IPPROTO_DIVERT (254)
value IPPROTO_DONE (257)
value IPPROTO_DSTOPTS (60)
value IPPROTO_EGP (8)
value IPPROTO_EMCON (14)
value IPPROTO_ENCAP (98)
value IPPROTO_EON (80)
value IPPROTO_ESP (50)
value IPPROTO_ETHERIP (97)
value IPPROTO_FRAGMENT (44)
value IPPROTO_GGP (3)
value IPPROTO_GMTP (100)
value IPPROTO_GRE (47)
value IPPROTO_HELLO (63)
value IPPROTO_HMP (20)
value IPPROTO_HOPOPTS (0)
value IPPROTO_ICMP (1)
value IPPROTO_IDP (22)
value IPPROTO_IDPR (35)
value IPPROTO_IDRP (45)
value IPPROTO_IGMP (2)
value IPPROTO_IGP (85)
value IPPROTO_IGRP (88)
value IPPROTO_IL (40)
value IPPROTO_INLSP (52)
value IPPROTO_INP (32)
value IPPROTO_IP (0)
value IPPROTO_IPCOMP (108)
value IPPROTO_IPCV (71)
value IPPROTO_IPEIP (94)
value IPPROTO_IPIP (IPPROTO_IPV4)
value IPPROTO_IPPC (67)
value IPPROTO_IRTP (28)
value IPPROTO_KRYPTOLAN (65)
value IPPROTO_LARP (91)
value IPPROTO_MAX (256)
value IPPROTO_MEAS (19)
value IPPROTO_MHRP (48)
value IPPROTO_MICP (95)
value IPPROTO_MTP (92)
value IPPROTO_MUX (18)
value IPPROTO_ND (77)
value IPPROTO_NHRP (54)
value IPPROTO_NONE (59)
value IPPROTO_NSP (31)
value IPPROTO_NVPII (11)
value IPPROTO_OSPFIGP (89)
value IPPROTO_PGM (113)
value IPPROTO_PIGP (9)
value IPPROTO_PIM (103)
value IPPROTO_PRM (21)
value IPPROTO_PUP (12)
value IPPROTO_PVP (75)
value IPPROTO_RAW (255)
value IPPROTO_RCCMON (10)
value IPPROTO_RDP (27)
value IPPROTO_ROUTING (43)
value IPPROTO_RSVP (46)
value IPPROTO_RVD (66)
value IPPROTO_SATEXPAK (64)
value IPPROTO_SATMON (69)
value IPPROTO_SCCSP (96)
value IPPROTO_SCTP (132)
value IPPROTO_SDRP (42)
value IPPROTO_SEP (33)
value IPPROTO_SRPC (90)
value IPPROTO_ST (7)
value IPPROTO_SVMTP (82)
value IPPROTO_SWIPE (53)
value IPPROTO_TCF (87)
value IPPROTO_TCP (6)
value IPPROTO_TP (29)
value IPPROTO_TPXX (39)
value IPPROTO_TTP (84)
value IPPROTO_UDP (17)
value IPPROTO_VINES (83)
value IPPROTO_VISA (70)
value IPPROTO_VMTP (81)
value IPPROTO_WBEXPAK (79)
value IPPROTO_WBMON (78)
value IPPROTO_WSN (74)
value IPPROTO_XNET (15)
value IPPROTO_XTP (36)
value IP_ADD_MEMBERSHIP (12)
value IP_ADD_SOURCE_MEMBERSHIP (70)
value IP_BLOCK_SOURCE (72)
value IP_BOUND_IF (25)
value IP_DEFAULT_MULTICAST_LOOP (1)
value IP_DEFAULT_MULTICAST_TTL (1)
value IP_DONTFRAG (28)
value IP_DROP_MEMBERSHIP (13)
value IP_DROP_SOURCE_MEMBERSHIP (71)
value IP_DUMMYNET_CONFIGURE (60)
value IP_DUMMYNET_DEL (61)
value IP_DUMMYNET_FLUSH (62)
value IP_DUMMYNET_GET (64)
value IP_FAITH (22)
value IP_FW_ADD (40)
value IP_FW_DEL (41)
value IP_FW_FLUSH (42)
value IP_FW_GET (44)
value IP_FW_RESETLOG (45)
value IP_FW_ZERO (43)
value IP_HDRINCL (2)
value IP_IPSEC_POLICY (21)
value IP_MAX_GROUP_SRC_FILTER (512)
value IP_MAX_MEMBERSHIPS (4095)
value IP_MAX_SOCK_MUTE_FILTER (128)
value IP_MAX_SOCK_SRC_FILTER (128)
value IP_MIN_MEMBERSHIPS (31)
value IP_MSFILTER (74)
value IP_MULTICAST_IF (9)
value IP_MULTICAST_IFINDEX (66)
value IP_MULTICAST_LOOP (11)
value IP_MULTICAST_TTL (10)
value IP_MULTICAST_VIF (14)
value IP_NAT__XXX (55)
value IP_OLD_FW_ADD (50)
value IP_OLD_FW_DEL (51)
value IP_OLD_FW_FLUSH (52)
value IP_OLD_FW_GET (54)
value IP_OLD_FW_RESETLOG (56)
value IP_OLD_FW_ZERO (53)
value IP_OPTIONS (1)
value IP_PKTINFO (26)
value IP_PORTRANGE (19)
value IP_PORTRANGE_DEFAULT (0)
value IP_PORTRANGE_HIGH (1)
value IP_PORTRANGE_LOW (2)
value IP_RECVDSTADDR (7)
value IP_RECVIF (20)
value IP_RECVOPTS (5)
value IP_RECVPKTINFO (IP_PKTINFO)
value IP_RECVRETOPTS (6)
value IP_RECVTOS (27)
value IP_RECVTTL (24)
value IP_RETOPTS (8)
value IP_RSVP_OFF (16)
value IP_RSVP_ON (15)
value IP_RSVP_VIF_OFF (18)
value IP_RSVP_VIF_ON (17)
value IP_STRIPHDR (23)
value IP_TOS (3)
value IP_TRAFFIC_MGT_BACKGROUND (65)
value IP_TTL (4)
value IP_UNBLOCK_SOURCE (73)
value ITIMER_PROF (2)
value ITIMER_REAL (0)
value ITIMER_VIRTUAL (1)
value KEV_DL_ADDMULTI (7)
value KEV_DL_AWDL_RESTRICTED (26)
value KEV_DL_AWDL_UNRESTRICTED (27)
value KEV_DL_DELMULTI (8)
value KEV_DL_IFCAP_CHANGED (19)
value KEV_DL_IFDELEGATE_CHANGED (25)
value KEV_DL_IF_ATTACHED (9)
value KEV_DL_IF_DETACHED (11)
value KEV_DL_IF_DETACHING (10)
value KEV_DL_IF_IDLE_ROUTE_REFCNT (18)
value KEV_DL_ISSUES (24)
value KEV_DL_LINK_ADDRESS_CHANGED (16)
value KEV_DL_LINK_OFF (12)
value KEV_DL_LINK_ON (13)
value KEV_DL_LINK_QUALITY_METRIC_CHANGED (20)
value KEV_DL_LOW_POWER_MODE_CHANGED (30)
value KEV_DL_MASTER_ELECTED (23)
value KEV_DL_NODE_ABSENCE (22)
value KEV_DL_NODE_PRESENCE (21)
value KEV_DL_PROTO_ATTACHED (14)
value KEV_DL_PROTO_DETACHED (15)
value KEV_DL_QOS_MODE_CHANGED (29)
value KEV_DL_RRC_STATE_CHANGED (28)
value KEV_DL_SIFFLAGS (1)
value KEV_DL_SIFGENERIC (6)
value KEV_DL_SIFMEDIA (5)
value KEV_DL_SIFMETRICS (2)
value KEV_DL_SIFMTU (3)
value KEV_DL_SIFPHYS (4)
value KEV_DL_SUBCLASS (2)
value KEV_DL_WAKEFLAGS_CHANGED (17)
value KEV_INET_ADDR_DELETED (3)
value KEV_INET_ARPCOLLISION (7)
value KEV_INET_ARPRTRALIVE (10)
value KEV_INET_ARPRTRFAILURE (9)
value KEV_INET_CHANGED_ADDR (2)
value KEV_INET_NEW_ADDR (1)
value KEV_INET_PORTINUSE (8)
value KEV_INET_SIFBRDADDR (5)
value KEV_INET_SIFDSTADDR (4)
value KEV_INET_SIFNETMASK (6)
value KEV_INET_SUBCLASS (1)
value LITTLE_ENDIAN (__DARWIN_LITTLE_ENDIAN)
value L_INCR (SEEK_CUR)
value L_SET (SEEK_SET)
value L_XTND (SEEK_END)
value MAXNAMLEN (__DARWIN_MAXNAMLEN)
value MCAST_BLOCK_SOURCE (84)
value MCAST_EXCLUDE (2)
value MCAST_INCLUDE (1)
value MCAST_JOIN_GROUP (80)
value MCAST_JOIN_SOURCE_GROUP (82)
value MCAST_LEAVE_GROUP (81)
value MCAST_LEAVE_SOURCE_GROUP (83)
value MCAST_UNBLOCK_SOURCE (85)
value MCAST_UNDEFINED (0)
value MINSIGSTKSZ (32768)
value NBBY (__DARWIN_NBBY)
value NETDB_SUCCESS (0)
value NETSVC_MRKNG_UNKNOWN (0)
value NET_MAXID (AF_MAX)
value NET_RT_DUMP (1)
value NET_RT_FLAGS (2)
value NET_RT_FLAGS_PRIV (10)
value NET_RT_IFLIST (3)
value NET_RT_MAXID (11)
value NET_RT_STAT (4)
value NET_RT_TRASH (5)
value NET_SERVICE_TYPE_AV (6)
value NET_SERVICE_TYPE_BE (0)
value NET_SERVICE_TYPE_BK (1)
value NET_SERVICE_TYPE_OAM (7)
value NET_SERVICE_TYPE_RD (8)
value NET_SERVICE_TYPE_RV (5)
value NET_SERVICE_TYPE_SIG (2)
value NET_SERVICE_TYPE_VI (3)
value NET_SERVICE_TYPE_VO (4)
value NFDBITS (__DARWIN_NFDBITS)
value NI_MAXHOST (1025)
value NI_MAXSERV (32)
value NO_ADDRESS (NO_DATA)
value NO_DATA (4)
value NO_RECOVERY (3)
value NSIG (__DARWIN_NSIG)
value NULL (__DARWIN_NULL)
value O_FSYNC (O_SYNC)
value O_NDELAY (O_NONBLOCK)
value PDP_ENDIAN (__DARWIN_PDP_ENDIAN)
value PF_APPLETALK (AF_APPLETALK)
value PF_CCITT (AF_CCITT)
value PF_CHAOS (AF_CHAOS)
value PF_CNT (AF_CNT)
value PF_COIP (AF_COIP)
value PF_DATAKIT (AF_DATAKIT)
value PF_DLI (AF_DLI)
value PF_ECMA (AF_ECMA)
value PF_HYLINK (AF_HYLINK)
value PF_IMPLINK (AF_IMPLINK)
value PF_INET (AF_INET)
value PF_IPX (AF_IPX)
value PF_ISDN (AF_ISDN)
value PF_ISO (AF_ISO)
value PF_LAT (AF_LAT)
value PF_LINK (AF_LINK)
value PF_LOCAL (AF_LOCAL)
value PF_MAX (AF_MAX)
value PF_NATM (AF_NATM)
value PF_NDRV (AF_NDRV)
value PF_NETBIOS (AF_NETBIOS)
value PF_NS (AF_NS)
value PF_OSI (AF_ISO)
value PF_PPP (AF_PPP)
value PF_PUP (AF_PUP)
value PF_ROUTE (AF_ROUTE)
value PF_SIP (AF_SIP)
value PF_SNA (AF_SNA)
value PF_SYSTEM (AF_SYSTEM)
value PF_UNIX (PF_LOCAL)
value PF_UNSPEC (AF_UNSPEC)
value PF_UTUN (AF_UTUN)
value PF_VSOCK (AF_VSOCK)
value POLLWRNORM (POLLOUT)
value POLL_ERR (4)
value POLL_HUP (6)
value POLL_IN (1)
value POLL_MSG (3)
value POLL_OUT (2)
value POLL_PRI (5)
value PRIO_DARWIN_PROCESS (4)
value PRIO_DARWIN_THREAD (3)
value PRIO_MAX (20)
value PRIO_PGRP (1)
value PRIO_PROCESS (0)
value PRIO_USER (2)
value PTRDIFF_MAX (INTMAX_MAX)
value PTRDIFF_MIN (INTMAX_MIN)
value RLIMIT_AS (5)
value RLIMIT_CORE (4)
value RLIMIT_CPU (0)
value RLIMIT_DATA (2)
value RLIMIT_FSIZE (1)
value RLIMIT_MEMLOCK (6)
value RLIMIT_NOFILE (8)
value RLIMIT_NPROC (7)
value RLIMIT_RSS (RLIMIT_AS)
value RLIMIT_STACK (3)
value RLIM_NLIMITS (9)
value RLIM_SAVED_CUR (RLIM_INFINITY)
value RLIM_SAVED_MAX (RLIM_INFINITY)
value RUSAGE_INFO_CURRENT (RUSAGE_INFO_V5)
value RUSAGE_SELF (0)
value SAE_ASSOCID_ANY (0)
value SAE_CONNID_ANY (0)
value SEEK_CUR (1)
value SEEK_DATA (4)
value SEEK_END (2)
value SEEK_HOLE (3)
value SEEK_SET (0)
value SEGV_ACCERR (2)
value SEGV_MAPERR (1)
value SEGV_NOOP (0)
value SHUT_RD (0)
value SHUT_RDWR (2)
value SHUT_WR (1)
value SIGABRT (6)
value SIGALRM (14)
value SIGBUS (10)
value SIGCHLD (20)
value SIGCONT (19)
value SIGEMT (7)
value SIGEV_NONE (0)
value SIGEV_SIGNAL (1)
value SIGEV_THREAD (3)
value SIGFPE (8)
value SIGHUP (1)
value SIGILL (4)
value SIGINFO (29)
value SIGINT (2)
value SIGIO (23)
value SIGIOT (SIGABRT)
value SIGKILL (9)
value SIGPIPE (13)
value SIGPROF (27)
value SIGQUIT (3)
value SIGSEGV (11)
value SIGSTKSZ (131072)
value SIGSTOP (17)
value SIGSYS (12)
value SIGTERM (15)
value SIGTRAP (5)
value SIGTSTP (18)
value SIGTTIN (21)
value SIGTTOU (22)
value SIGURG (16)
value SIGVTALRM (26)
value SIGWINCH (28)
value SIGXCPU (24)
value SIGXFSZ (25)
value SIG_ATOMIC_MAX (INT32_MAX)
value SIG_ATOMIC_MIN (INT32_MIN)
value SIG_BLOCK (1)
value SIG_SETMASK (3)
value SIG_UNBLOCK (2)
value SIZE_MAX (UINTPTR_MAX)
value SOCK_DGRAM (2)
value SOCK_MAXADDRLEN (255)
value SOCK_RAW (3)
value SOCK_RDM (4)
value SOCK_SEQPACKET (5)
value SOCK_STREAM (1)
value SOMAXCONN (128)
value STDERR_FILENO (2)
value STDIN_FILENO (0)
value STDOUT_FILENO (1)
value SV_INTERRUPT (SA_RESTART)
value SV_NOCLDSTOP (SA_NOCLDSTOP)
value SV_NODEFER (SA_NODEFER)
value SV_ONSTACK (SA_ONSTACK)
value SV_RESETHAND (SA_RESETHAND)
value SV_SIGINFO (SA_SIGINFO)
value S_BLKSIZE (512)
value S_IEXEC (S_IXUSR)
value S_IFBLK (0c060000)
value S_IFCHR (0c020000)
value S_IFDIR (0c040000)
value S_IFIFO (0c010000)
value S_IFLNK (0c120000)
value S_IFMT (0c170000)
value S_IFREG (0c100000)
value S_IFSOCK (0c140000)
value S_IFWHT (0c160000)
value S_IREAD (S_IRUSR)
value S_IRGRP (0c000040)
value S_IROTH (0c000004)
value S_IRUSR (0c000400)
value S_IRWXG (0c000070)
value S_IRWXO (0c000007)
value S_IRWXU (0c000700)
value S_ISGID (0c002000)
value S_ISTXT (S_ISVTX)
value S_ISUID (0c004000)
value S_ISVTX (0c001000)
value S_IWGRP (0c000020)
value S_IWOTH (0c000002)
value S_IWRITE (S_IWUSR)
value S_IWUSR (0c000200)
value S_IXGRP (0c000010)
value S_IXOTH (0c000001)
value S_IXUSR (0c000100)
value TIME_UTC (1)
value TMP_MAX (308915776)
value TRAP_BRKPT (1)
value TRAP_TRACE (2)
value TRY_AGAIN (2)
value UINTPTR_MAX (18446744073709551615UL)
value USER_FSIGNATURES_CDHASH_LEN (20)
value WAIT_MYPGRP (0)
value WCHAR_MAX (__WCHAR_MAX__)
value WCOREFLAG (0c200)
value WINT_MAX (INT32_MAX)
value WINT_MIN (INT32_MIN)
value _ARM_SIGNAL_ (1)
value _CS_DARWIN_USER_CACHE_DIR (65538)
value _CS_DARWIN_USER_DIR (65536)
value _CS_DARWIN_USER_TEMP_DIR (65537)
value _CS_PATH (1)
value _DARWIN_FEATURE_ONLY_UNIX_CONFORMANCE (1)
value _DARWIN_FEATURE_UNIX_CONFORMANCE (3)
value _FORTIFY_SOURCE (0)
value _IOFBF (0)
value _IOLBF (1)
value _IONBF (2)
value _PC_ALLOC_SIZE_MIN (16)
value _PC_ASYNC_IO (17)
value _PC_AUTH_OPAQUE_NP (14)
value _PC_CASE_PRESERVING (12)
value _PC_CASE_SENSITIVE (11)
value _PC_CHOWN_RESTRICTED (7)
value _PC_EXTENDED_SECURITY_NP (13)
value _PC_FILESIZEBITS (18)
value _PC_LINK_MAX (1)
value _PC_MAX_CANON (2)
value _PC_MAX_INPUT (3)
value _PC_MIN_HOLE_SIZE (27)
value _PC_NAME_CHARS_MAX (10)
value _PC_NAME_MAX (4)
value _PC_NO_TRUNC (8)
value _PC_PATH_MAX (5)
value _PC_PIPE_BUF (6)
value _PC_PRIO_IO (19)
value _PC_REC_INCR_XFER_SIZE (20)
value _PC_REC_MAX_XFER_SIZE (21)
value _PC_REC_MIN_XFER_SIZE (22)
value _PC_REC_XFER_ALIGN (23)
value _PC_SYMLINK_MAX (24)
value _PC_SYNC_IO (25)
value _PC_VDISABLE (9)
value _PC_XATTR_SIZE_BITS (26)
value _POSIX_CHOWN_RESTRICTED (200112L)
value _POSIX_FSYNC (200112L)
value _POSIX_JOB_CONTROL (200112L)
value _POSIX_MAPPED_FILES (200112L)
value _POSIX_MEMORY_PROTECTION (200112L)
value _POSIX_NO_TRUNC (200112L)
value _POSIX_READER_WRITER_LOCKS (200112L)
value _POSIX_REGEXP (200112L)
value _POSIX_SAVED_IDS (200112L)
value _POSIX_SHELL (200112L)
value _POSIX_THREADS (200112L)
value _POSIX_THREAD_ATTR_STACKADDR (200112L)
value _POSIX_THREAD_ATTR_STACKSIZE (200112L)
value _POSIX_THREAD_KEYS_MAX (128)
value _POSIX_THREAD_PROCESS_SHARED (200112L)
value _POSIX_THREAD_SAFE_FUNCTIONS (200112L)
value _POSIX_VERSION (200112L)
value _QUAD_HIGHWORD (1)
value _QUAD_LOWWORD (0)
value _SC_ADVISORY_INFO (65)
value _SC_AIO_LISTIO_MAX (42)
value _SC_AIO_MAX (43)
value _SC_AIO_PRIO_DELTA_MAX (44)
value _SC_ARG_MAX (1)
value _SC_ASYNCHRONOUS_IO (28)
value _SC_ATEXIT_MAX (107)
value _SC_BARRIERS (66)
value _SC_BC_BASE_MAX (9)
value _SC_BC_DIM_MAX (10)
value _SC_BC_SCALE_MAX (11)
value _SC_BC_STRING_MAX (12)
value _SC_CHILD_MAX (2)
value _SC_CLK_TCK (3)
value _SC_CLOCK_SELECTION (67)
value _SC_COLL_WEIGHTS_MAX (13)
value _SC_CPUTIME (68)
value _SC_DELAYTIMER_MAX (45)
value _SC_EXPR_NEST_MAX (14)
value _SC_FILE_LOCKING (69)
value _SC_FSYNC (38)
value _SC_GETGR_R_SIZE_MAX (70)
value _SC_GETPW_R_SIZE_MAX (71)
value _SC_HOST_NAME_MAX (72)
value _SC_IOV_MAX (56)
value _SC_JOB_CONTROL (6)
value _SC_LINE_MAX (15)
value _SC_LOGIN_NAME_MAX (73)
value _SC_MAPPED_FILES (47)
value _SC_MEMLOCK (30)
value _SC_MEMLOCK_RANGE (31)
value _SC_MEMORY_PROTECTION (32)
value _SC_MESSAGE_PASSING (33)
value _SC_MONOTONIC_CLOCK (74)
value _SC_MQ_OPEN_MAX (46)
value _SC_MQ_PRIO_MAX (75)
value _SC_NGROUPS_MAX (4)
value _SC_NPROCESSORS_CONF (57)
value _SC_NPROCESSORS_ONLN (58)
value _SC_OPEN_MAX (5)
value _SC_PAGESIZE (29)
value _SC_PAGE_SIZE (_SC_PAGESIZE)
value _SC_PASS_MAX (131)
value _SC_PHYS_PAGES (200)
value _SC_PRIORITIZED_IO (34)
value _SC_PRIORITY_SCHEDULING (35)
value _SC_RAW_SOCKETS (119)
value _SC_READER_WRITER_LOCKS (76)
value _SC_REALTIME_SIGNALS (36)
value _SC_REGEXP (77)
value _SC_RE_DUP_MAX (16)
value _SC_RTSIG_MAX (48)
value _SC_SAVED_IDS (7)
value _SC_SEMAPHORES (37)
value _SC_SEM_NSEMS_MAX (49)
value _SC_SEM_VALUE_MAX (50)
value _SC_SHARED_MEMORY_OBJECTS (39)
value _SC_SHELL (78)
value _SC_SIGQUEUE_MAX (51)
value _SC_SPAWN (79)
value _SC_SPIN_LOCKS (80)
value _SC_SPORADIC_SERVER (81)
value _SC_SS_REPL_MAX (126)
value _SC_STREAM_MAX (26)
value _SC_SYMLOOP_MAX (120)
value _SC_SYNCHRONIZED_IO (40)
value _SC_THREADS (96)
value _SC_THREAD_ATTR_STACKADDR (82)
value _SC_THREAD_ATTR_STACKSIZE (83)
value _SC_THREAD_CPUTIME (84)
value _SC_THREAD_DESTRUCTOR_ITERATIONS (85)
value _SC_THREAD_KEYS_MAX (86)
value _SC_THREAD_PRIORITY_SCHEDULING (89)
value _SC_THREAD_PRIO_INHERIT (87)
value _SC_THREAD_PRIO_PROTECT (88)
value _SC_THREAD_PROCESS_SHARED (90)
value _SC_THREAD_SAFE_FUNCTIONS (91)
value _SC_THREAD_SPORADIC_SERVER (92)
value _SC_THREAD_STACK_MIN (93)
value _SC_THREAD_THREADS_MAX (94)
value _SC_TIMEOUTS (95)
value _SC_TIMERS (41)
value _SC_TIMER_MAX (52)
value _SC_TRACE (97)
value _SC_TRACE_EVENT_FILTER (98)
value _SC_TRACE_EVENT_NAME_MAX (127)
value _SC_TRACE_INHERIT (99)
value _SC_TRACE_LOG (100)
value _SC_TRACE_NAME_MAX (128)
value _SC_TRACE_SYS_MAX (129)
value _SC_TRACE_USER_EVENT_MAX (130)
value _SC_TTY_NAME_MAX (101)
value _SC_TYPED_MEMORY_OBJECTS (102)
value _SC_TZNAME_MAX (27)
value _SC_VERSION (8)
value _SC_XOPEN_CRYPT (108)
value _SC_XOPEN_LEGACY (110)
value _SC_XOPEN_REALTIME (111)
value _SC_XOPEN_REALTIME_THREADS (112)
value _SC_XOPEN_SHM (113)
value _SC_XOPEN_STREAMS (114)
value _SC_XOPEN_UNIX (115)
value _SC_XOPEN_VERSION (116)
value _SC_XOPEN_XCU_VERSION (121)
value _SS_MAXSIZE (128)
value _STRUCT_MCONTEXT (_STRUCT_MCONTEXT64)
value _WSTOPPED (0c177)
value _XOPEN_VERSION (600)
value _XOPEN_XCU_VERSION (4)
value __API_TO_BE_DEPRECATED (100000)
value __APPLE_CC__ (6000)
value __APPLE__ (1)
value __ARM_ACLE (200)
value __ARM_ALIGN_MAX_STACK_PWR (4)
value __ARM_ARCH (8)
value __ARM_FEATURE_AES (1)
value __ARM_FEATURE_ATOMICS (1)
value __ARM_FEATURE_CLZ (1)
value __ARM_FEATURE_COMPLEX (1)
value __ARM_FEATURE_CRYPTO (1)
value __ARM_FEATURE_DIRECTED_ROUNDING (1)
value __ARM_FEATURE_DIV (1)
value __ARM_FEATURE_DOTPROD (1)
value __ARM_FEATURE_FMA (1)
value __ARM_FEATURE_FRINT (1)
value __ARM_FEATURE_IDIV (1)
value __ARM_FEATURE_JCVT (1)
value __ARM_FEATURE_NUMERIC_MAXMIN (1)
value __ARM_FEATURE_QRDMX (1)
value __ARM_FEATURE_UNALIGNED (1)
value __ARM_NEON (1)
value __ARM_NEON__ (1)
value __ARM_SIZEOF_MINIMAL_ENUM (4)
value __ARM_SIZEOF_WCHAR_T (4)
value __ATOMIC_ACQUIRE (2)
value __ATOMIC_ACQ_REL (4)
value __ATOMIC_CONSUME (1)
value __ATOMIC_RELAXED (0)
value __ATOMIC_RELEASE (3)
value __ATOMIC_SEQ_CST (5)
value __BIGGEST_ALIGNMENT__ (8)
value __BITINT_MAXWIDTH__ (128)
value __BLOCKS__ (1)
value __BOOL_WIDTH__ (8)
value __BYTE_ORDER__ (__ORDER_LITTLE_ENDIAN__)
value __CHAR_BIT__ (8)
value __CLANG_ATOMIC_BOOL_LOCK_FREE (2)
value __CLANG_ATOMIC_CHAR_LOCK_FREE (2)
value __CLANG_ATOMIC_INT_LOCK_FREE (2)
value __CLANG_ATOMIC_LLONG_LOCK_FREE (2)
value __CLANG_ATOMIC_LONG_LOCK_FREE (2)
value __CLANG_ATOMIC_POINTER_LOCK_FREE (2)
value __CLANG_ATOMIC_SHORT_LOCK_FREE (2)
value __CLANG_ATOMIC_WCHAR_T_LOCK_FREE (2)
value __CONSTANT_CFSTRINGS__ (1)
value __DARWIN_BIG_ENDIAN (4321)
value __DARWIN_BYTE_ORDER (__DARWIN_LITTLE_ENDIAN)
value __DARWIN_C_ANSI (0c10000L)
value __DARWIN_C_FULL (900000L)
value __DARWIN_C_LEVEL (__DARWIN_C_FULL)
value __DARWIN_FD_SETSIZE (1024)
value __DARWIN_IPPORT_RESERVED (1024)
value __DARWIN_LITTLE_ENDIAN (1234)
value __DARWIN_MAXNAMLEN (255)
value __DARWIN_MAXPATHLEN (1024)
value __DARWIN_NBBY (8)
value __DARWIN_NON_CANCELABLE (0)
value __DARWIN_NO_LONG_LONG (0)
value __DARWIN_NSIG (32)
value __DARWIN_ONLY_UNIX_CONFORMANCE (1)
value __DARWIN_PDP_ENDIAN (3412)
value __DARWIN_WCHAR_MAX (__WCHAR_MAX__)
value __DBL_DECIMAL_DIG__ (17)
value __DBL_DIG__ (15)
value __DBL_HAS_DENORM__ (1)
value __DBL_HAS_INFINITY__ (1)
value __DBL_HAS_QUIET_NAN__ (1)
value __DBL_MANT_DIG__ (53)
value __DBL_MAX_EXP__ (1024)
value __DECIMAL_DIG__ (__LDBL_DECIMAL_DIG__)
value __DYNAMIC__ (1)
value __ENABLE_LEGACY_MAC_AVAILABILITY (1)
value __ENVIRONMENT_MAC_OS_X_VERSION_MIN_REQUIRED__ (1040)
value __FINITE_MATH_ONLY__ (0)
value __FLT_DECIMAL_DIG__ (9)
value __FLT_DIG__ (6)
value __FLT_HAS_DENORM__ (1)
value __FLT_HAS_INFINITY__ (1)
value __FLT_HAS_QUIET_NAN__ (1)
value __FLT_MANT_DIG__ (24)
value __FLT_MAX_EXP__ (128)
value __FLT_RADIX__ (2)
value __FP_FAST_FMA (1)
value __FP_FAST_FMAF (1)
value __GCC_ATOMIC_BOOL_LOCK_FREE (2)
value __GCC_ATOMIC_CHAR_LOCK_FREE (2)
value __GCC_ATOMIC_INT_LOCK_FREE (2)
value __GCC_ATOMIC_LLONG_LOCK_FREE (2)
value __GCC_ATOMIC_LONG_LOCK_FREE (2)
value __GCC_ATOMIC_POINTER_LOCK_FREE (2)
value __GCC_ATOMIC_SHORT_LOCK_FREE (2)
value __GCC_ATOMIC_TEST_AND_SET_TRUEVAL (1)
value __GCC_ATOMIC_WCHAR_T_LOCK_FREE (2)
value __GNUC_MINOR__ (2)
value __GNUC_PATCHLEVEL__ (1)
value __GNUC_STDC_INLINE__ (1)
value __GNUC__ (4)
value __GXX_ABI_VERSION (1002)
value __INTMAX_C_SUFFIX__ (L)
value __INTMAX_MAX__ (9223372036854775807L)
value __INTMAX_WIDTH__ (64)
value __INTPTR_MAX__ (9223372036854775807L)
value __INTPTR_WIDTH__ (64)
value __INT_MAX__ (2147483647)
value __INT_WIDTH__ (32)
value __LDBL_DECIMAL_DIG__ (17)
value __LDBL_DIG__ (15)
value __LDBL_HAS_DENORM__ (1)
value __LDBL_HAS_INFINITY__ (1)
value __LDBL_HAS_QUIET_NAN__ (1)
value __LDBL_MANT_DIG__ (53)
value __LDBL_MAX_EXP__ (1024)
value __LITTLE_ENDIAN__ (1)
value __LLONG_WIDTH__ (64)
value __LONG_LONG_MAX__ (9223372036854775807LL)
value __LONG_MAX__ (9223372036854775807L)
value __LONG_WIDTH__ (64)
value __MACH__ (1)
value __MAC_OS_X_VERSION_MAX_ALLOWED (__MAC_11_3)
value __MAC_OS_X_VERSION_MIN_REQUIRED (__ENVIRONMENT_MAC_OS_X_VERSION_MIN_REQUIRED__)
value __NO_INLINE__ (1)
value __NO_MATH_ERRNO__ (1)
value __OBJC_BOOL_IS_BOOL (1)
value __OPENCL_MEMORY_SCOPE_ALL_SVM_DEVICES (3)
value __OPENCL_MEMORY_SCOPE_DEVICE (2)
value __OPENCL_MEMORY_SCOPE_SUB_GROUP (4)
value __OPENCL_MEMORY_SCOPE_WORK_GROUP (1)
value __OPENCL_MEMORY_SCOPE_WORK_ITEM (0)
value __ORDER_BIG_ENDIAN__ (4321)
value __ORDER_LITTLE_ENDIAN__ (1234)
value __ORDER_PDP_ENDIAN__ (3412)
value __PIC__ (2)
value __POINTER_WIDTH__ (64)
value __PRAGMA_REDEFINE_EXTNAME (1)
value __PTHREAD_ATTR_SIZE__ (56)
value __PTHREAD_CONDATTR_SIZE__ (8)
value __PTHREAD_COND_SIZE__ (40)
value __PTHREAD_MUTEXATTR_SIZE__ (8)
value __PTHREAD_MUTEX_SIZE__ (56)
value __PTHREAD_ONCE_SIZE__ (8)
value __PTHREAD_RWLOCKATTR_SIZE__ (16)
value __PTHREAD_RWLOCK_SIZE__ (192)
value __PTHREAD_SIZE__ (8176)
value __PTRDIFF_MAX__ (9223372036854775807L)
value __PTRDIFF_WIDTH__ (64)
value __SCHAR_MAX__ (127)
value __SHRT_MAX__ (32767)
value __SHRT_WIDTH__ (16)
value __SIG_ATOMIC_MAX__ (2147483647)
value __SIG_ATOMIC_WIDTH__ (32)
value __SIZEOF_DOUBLE__ (8)
value __SIZEOF_FLOAT__ (4)
value __SIZEOF_INT__ (4)
value __SIZEOF_LONG_DOUBLE__ (8)
value __SIZEOF_LONG_LONG__ (8)
value __SIZEOF_LONG__ (8)
value __SIZEOF_POINTER__ (8)
value __SIZEOF_PTRDIFF_T__ (8)
value __SIZEOF_SHORT__ (2)
value __SIZEOF_SIZE_T__ (8)
value __SIZEOF_WCHAR_T__ (4)
value __SIZEOF_WINT_T__ (4)
value __SIZE_MAX__ (18446744073709551615UL)
value __SIZE_WIDTH__ (64)
value __SSP__ (1)
value __STDC_HOSTED__ (1)
value __STDC_NO_THREADS__ (1)
value __STDC_VERSION__ (201710L)
value __STDC__ (1)
value __UINTMAX_C_SUFFIX__ (UL)
value __UINTMAX_MAX__ (18446744073709551615UL)
value __UINTMAX_WIDTH__ (64)
value __UINTPTR_MAX__ (18446744073709551615UL)
value __UINTPTR_WIDTH__ (64)
value __USER_LABEL_PREFIX__ (_)
value __WCHAR_MAX__ (2147483647)
value __WCHAR_WIDTH__ (32)
value __WINT_MAX__ (2147483647)
value __WINT_WIDTH__ (32)
value __WORDSIZE (64)

